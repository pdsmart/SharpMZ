-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b83ff",
             1 => x"f80d0b0b",
             2 => x"0b93b904",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"9d040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b9380",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b8295",
           162 => x"bc738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93850400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b80c3",
           171 => x"f42d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b80c5",
           179 => x"e02d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"95040b0b",
           269 => x"0b8ca404",
           270 => x"0b0b0b8c",
           271 => x"b3040b0b",
           272 => x"0b8cc204",
           273 => x"0b0b0b8c",
           274 => x"d1040b0b",
           275 => x"0b8ce004",
           276 => x"0b0b0b8c",
           277 => x"f0040b0b",
           278 => x"0b8d8004",
           279 => x"0b0b0b8d",
           280 => x"8f040b0b",
           281 => x"0b8d9e04",
           282 => x"0b0b0b8d",
           283 => x"ad040b0b",
           284 => x"0b8dbd04",
           285 => x"0b0b0b8d",
           286 => x"cd040b0b",
           287 => x"0b8ddd04",
           288 => x"0b0b0b8d",
           289 => x"ed040b0b",
           290 => x"0b8dfd04",
           291 => x"0b0b0b8e",
           292 => x"8d040b0b",
           293 => x"0b8e9d04",
           294 => x"0b0b0b8e",
           295 => x"ad040b0b",
           296 => x"0b8ebd04",
           297 => x"0b0b0b8e",
           298 => x"cd040b0b",
           299 => x"0b8edd04",
           300 => x"0b0b0b8e",
           301 => x"ed040b0b",
           302 => x"0b8efd04",
           303 => x"0b0b0b8f",
           304 => x"8d040b0b",
           305 => x"0b8f9d04",
           306 => x"0b0b0b8f",
           307 => x"ad040b0b",
           308 => x"0b8fbd04",
           309 => x"0b0b0b8f",
           310 => x"cd040b0b",
           311 => x"0b8fdd04",
           312 => x"0b0b0b8f",
           313 => x"ed040b0b",
           314 => x"0b8ffd04",
           315 => x"0b0b0b90",
           316 => x"8d040b0b",
           317 => x"0b909d04",
           318 => x"0b0b0b90",
           319 => x"ad040b0b",
           320 => x"0b90bd04",
           321 => x"0b0b0b90",
           322 => x"cd040b0b",
           323 => x"0b90dd04",
           324 => x"0b0b0b90",
           325 => x"ed040b0b",
           326 => x"0b90fd04",
           327 => x"0b0b0b91",
           328 => x"8d040b0b",
           329 => x"0b919d04",
           330 => x"0b0b0b91",
           331 => x"ad040b0b",
           332 => x"0b91bd04",
           333 => x"0b0b0b91",
           334 => x"cd040b0b",
           335 => x"0b91dd04",
           336 => x"0b0b0b91",
           337 => x"ed040b0b",
           338 => x"0b91fd04",
           339 => x"0b0b0b92",
           340 => x"8d040b0b",
           341 => x"0b929d04",
           342 => x"0b0b0b92",
           343 => x"ad040b0b",
           344 => x"0b92bd04",
           345 => x"0b0b0b92",
           346 => x"cd04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0482b6a4",
           386 => x"0c80f4fe",
           387 => x"2d82b6a4",
           388 => x"0882d090",
           389 => x"0482b6a4",
           390 => x"0cb3b22d",
           391 => x"82b6a408",
           392 => x"82d09004",
           393 => x"82b6a40c",
           394 => x"afe32d82",
           395 => x"b6a40882",
           396 => x"d0900482",
           397 => x"b6a40caf",
           398 => x"ad2d82b6",
           399 => x"a40882d0",
           400 => x"900482b6",
           401 => x"a40c94ad",
           402 => x"2d82b6a4",
           403 => x"0882d090",
           404 => x"0482b6a4",
           405 => x"0cb1c22d",
           406 => x"82b6a408",
           407 => x"82d09004",
           408 => x"82b6a40c",
           409 => x"80cfcc2d",
           410 => x"82b6a408",
           411 => x"82d09004",
           412 => x"82b6a40c",
           413 => x"80c9fb2d",
           414 => x"82b6a408",
           415 => x"82d09004",
           416 => x"82b6a40c",
           417 => x"93d82d82",
           418 => x"b6a40882",
           419 => x"d0900482",
           420 => x"b6a40c96",
           421 => x"c02d82b6",
           422 => x"a40882d0",
           423 => x"900482b6",
           424 => x"a40c97cd",
           425 => x"2d82b6a4",
           426 => x"0882d090",
           427 => x"0482b6a4",
           428 => x"0c80f8a8",
           429 => x"2d82b6a4",
           430 => x"0882d090",
           431 => x"0482b6a4",
           432 => x"0c80f986",
           433 => x"2d82b6a4",
           434 => x"0882d090",
           435 => x"0482b6a4",
           436 => x"0c80f0c3",
           437 => x"2d82b6a4",
           438 => x"0882d090",
           439 => x"0482b6a4",
           440 => x"0c80f2ba",
           441 => x"2d82b6a4",
           442 => x"0882d090",
           443 => x"0482b6a4",
           444 => x"0c80f3ed",
           445 => x"2d82b6a4",
           446 => x"0882d090",
           447 => x"0482b6a4",
           448 => x"0c81d89e",
           449 => x"2d82b6a4",
           450 => x"0882d090",
           451 => x"0482b6a4",
           452 => x"0c81e58f",
           453 => x"2d82b6a4",
           454 => x"0882d090",
           455 => x"0482b6a4",
           456 => x"0c81dd83",
           457 => x"2d82b6a4",
           458 => x"0882d090",
           459 => x"0482b6a4",
           460 => x"0c81e080",
           461 => x"2d82b6a4",
           462 => x"0882d090",
           463 => x"0482b6a4",
           464 => x"0c81ea9e",
           465 => x"2d82b6a4",
           466 => x"0882d090",
           467 => x"0482b6a4",
           468 => x"0c81f2fe",
           469 => x"2d82b6a4",
           470 => x"0882d090",
           471 => x"0482b6a4",
           472 => x"0c81e3f1",
           473 => x"2d82b6a4",
           474 => x"0882d090",
           475 => x"0482b6a4",
           476 => x"0c81edbd",
           477 => x"2d82b6a4",
           478 => x"0882d090",
           479 => x"0482b6a4",
           480 => x"0c81eedc",
           481 => x"2d82b6a4",
           482 => x"0882d090",
           483 => x"0482b6a4",
           484 => x"0c81eefb",
           485 => x"2d82b6a4",
           486 => x"0882d090",
           487 => x"0482b6a4",
           488 => x"0c81f6e5",
           489 => x"2d82b6a4",
           490 => x"0882d090",
           491 => x"0482b6a4",
           492 => x"0c81f4cb",
           493 => x"2d82b6a4",
           494 => x"0882d090",
           495 => x"0482b6a4",
           496 => x"0c81f9b9",
           497 => x"2d82b6a4",
           498 => x"0882d090",
           499 => x"0482b6a4",
           500 => x"0c81efff",
           501 => x"2d82b6a4",
           502 => x"0882d090",
           503 => x"0482b6a4",
           504 => x"0c81fcb9",
           505 => x"2d82b6a4",
           506 => x"0882d090",
           507 => x"0482b6a4",
           508 => x"0c81fdba",
           509 => x"2d82b6a4",
           510 => x"0882d090",
           511 => x"0482b6a4",
           512 => x"0c81e5ef",
           513 => x"2d82b6a4",
           514 => x"0882d090",
           515 => x"0482b6a4",
           516 => x"0c81e5c8",
           517 => x"2d82b6a4",
           518 => x"0882d090",
           519 => x"0482b6a4",
           520 => x"0c81e6f3",
           521 => x"2d82b6a4",
           522 => x"0882d090",
           523 => x"0482b6a4",
           524 => x"0c81f0d6",
           525 => x"2d82b6a4",
           526 => x"0882d090",
           527 => x"0482b6a4",
           528 => x"0c81feab",
           529 => x"2d82b6a4",
           530 => x"0882d090",
           531 => x"0482b6a4",
           532 => x"0c8280b5",
           533 => x"2d82b6a4",
           534 => x"0882d090",
           535 => x"0482b6a4",
           536 => x"0c8283f7",
           537 => x"2d82b6a4",
           538 => x"0882d090",
           539 => x"0482b6a4",
           540 => x"0c81d7bd",
           541 => x"2d82b6a4",
           542 => x"0882d090",
           543 => x"0482b6a4",
           544 => x"0c8286e3",
           545 => x"2d82b6a4",
           546 => x"0882d090",
           547 => x"0482b6a4",
           548 => x"0c829598",
           549 => x"2d82b6a4",
           550 => x"0882d090",
           551 => x"0482b6a4",
           552 => x"0c829384",
           553 => x"2d82b6a4",
           554 => x"0882d090",
           555 => x"0482b6a4",
           556 => x"0c81a8f8",
           557 => x"2d82b6a4",
           558 => x"0882d090",
           559 => x"0482b6a4",
           560 => x"0c81aae2",
           561 => x"2d82b6a4",
           562 => x"0882d090",
           563 => x"0482b6a4",
           564 => x"0c81acc6",
           565 => x"2d82b6a4",
           566 => x"0882d090",
           567 => x"0482b6a4",
           568 => x"0c80f0ec",
           569 => x"2d82b6a4",
           570 => x"0882d090",
           571 => x"0482b6a4",
           572 => x"0c80f290",
           573 => x"2d82b6a4",
           574 => x"0882d090",
           575 => x"0482b6a4",
           576 => x"0c80f5f3",
           577 => x"2d82b6a4",
           578 => x"0882d090",
           579 => x"0482b6a4",
           580 => x"0c80d698",
           581 => x"2d82b6a4",
           582 => x"0882d090",
           583 => x"0482b6a4",
           584 => x"0c81a38c",
           585 => x"2d82b6a4",
           586 => x"0882d090",
           587 => x"0482b6a4",
           588 => x"0c81a3b4",
           589 => x"2d82b6a4",
           590 => x"0882d090",
           591 => x"0482b6a4",
           592 => x"0c81a7ac",
           593 => x"2d82b6a4",
           594 => x"0882d090",
           595 => x"0482b6a4",
           596 => x"0c819ff6",
           597 => x"2d82b6a4",
           598 => x"0882d090",
           599 => x"043c0400",
           600 => x"00101010",
           601 => x"10101010",
           602 => x"10101010",
           603 => x"10101010",
           604 => x"10101010",
           605 => x"10101010",
           606 => x"10101010",
           607 => x"10101010",
           608 => x"53510400",
           609 => x"007381ff",
           610 => x"06738306",
           611 => x"09810583",
           612 => x"05101010",
           613 => x"2b0772fc",
           614 => x"060c5151",
           615 => x"04727280",
           616 => x"728106ff",
           617 => x"05097206",
           618 => x"05711052",
           619 => x"720a100a",
           620 => x"5372ed38",
           621 => x"51515351",
           622 => x"0482b698",
           623 => x"7082cdf4",
           624 => x"278e3880",
           625 => x"71708405",
           626 => x"530c0b0b",
           627 => x"0b93bc04",
           628 => x"8c815180",
           629 => x"ef860400",
           630 => x"82b6a408",
           631 => x"0282b6a4",
           632 => x"0cfb3d0d",
           633 => x"82b6a408",
           634 => x"8c057082",
           635 => x"b6a408fc",
           636 => x"050c82b6",
           637 => x"a408fc05",
           638 => x"085482b6",
           639 => x"a4088805",
           640 => x"085382cd",
           641 => x"ec085254",
           642 => x"849a3f82",
           643 => x"b6980870",
           644 => x"82b6a408",
           645 => x"f8050c82",
           646 => x"b6a408f8",
           647 => x"05087082",
           648 => x"b6980c51",
           649 => x"54873d0d",
           650 => x"82b6a40c",
           651 => x"0482b6a4",
           652 => x"080282b6",
           653 => x"a40cfb3d",
           654 => x"0d82b6a4",
           655 => x"08900508",
           656 => x"85113370",
           657 => x"81327081",
           658 => x"06515151",
           659 => x"52718f38",
           660 => x"800b82b6",
           661 => x"a4088c05",
           662 => x"08258338",
           663 => x"8d39800b",
           664 => x"82b6a408",
           665 => x"f4050c81",
           666 => x"c43982b6",
           667 => x"a4088c05",
           668 => x"08ff0582",
           669 => x"b6a4088c",
           670 => x"050c800b",
           671 => x"82b6a408",
           672 => x"f8050c82",
           673 => x"b6a40888",
           674 => x"050882b6",
           675 => x"a408fc05",
           676 => x"0c82b6a4",
           677 => x"08f80508",
           678 => x"8a2e80f6",
           679 => x"38800b82",
           680 => x"b6a4088c",
           681 => x"05082580",
           682 => x"e93882b6",
           683 => x"a4089005",
           684 => x"0851a090",
           685 => x"3f82b698",
           686 => x"087082b6",
           687 => x"a408f805",
           688 => x"0c5282b6",
           689 => x"a408f805",
           690 => x"08ff2e09",
           691 => x"81068d38",
           692 => x"800b82b6",
           693 => x"a408f405",
           694 => x"0c80d239",
           695 => x"82b6a408",
           696 => x"fc050882",
           697 => x"b6a408f8",
           698 => x"05085353",
           699 => x"71733482",
           700 => x"b6a4088c",
           701 => x"0508ff05",
           702 => x"82b6a408",
           703 => x"8c050c82",
           704 => x"b6a408fc",
           705 => x"05088105",
           706 => x"82b6a408",
           707 => x"fc050cff",
           708 => x"803982b6",
           709 => x"a408fc05",
           710 => x"08528072",
           711 => x"3482b6a4",
           712 => x"08880508",
           713 => x"7082b6a4",
           714 => x"08f4050c",
           715 => x"5282b6a4",
           716 => x"08f40508",
           717 => x"82b6980c",
           718 => x"873d0d82",
           719 => x"b6a40c04",
           720 => x"82b6a408",
           721 => x"0282b6a4",
           722 => x"0cf43d0d",
           723 => x"860b82b6",
           724 => x"a408e505",
           725 => x"3482b6a4",
           726 => x"08880508",
           727 => x"82b6a408",
           728 => x"e0050cfe",
           729 => x"0a0b82b6",
           730 => x"a408e805",
           731 => x"0c82b6a4",
           732 => x"08900570",
           733 => x"82b6a408",
           734 => x"fc050c82",
           735 => x"b6a408fc",
           736 => x"05085482",
           737 => x"b6a4088c",
           738 => x"05085382",
           739 => x"b6a408e0",
           740 => x"05705351",
           741 => x"54818d3f",
           742 => x"82b69808",
           743 => x"7082b6a4",
           744 => x"08dc050c",
           745 => x"82b6a408",
           746 => x"ec050882",
           747 => x"b6a40888",
           748 => x"05080551",
           749 => x"54807434",
           750 => x"82b6a408",
           751 => x"dc050870",
           752 => x"82b6980c",
           753 => x"548e3d0d",
           754 => x"82b6a40c",
           755 => x"0482b6a4",
           756 => x"080282b6",
           757 => x"a40cfb3d",
           758 => x"0d82b6a4",
           759 => x"08900570",
           760 => x"82b6a408",
           761 => x"fc050c82",
           762 => x"b6a408fc",
           763 => x"05085482",
           764 => x"b6a4088c",
           765 => x"05085382",
           766 => x"b6a40888",
           767 => x"05085254",
           768 => x"a33f82b6",
           769 => x"98087082",
           770 => x"b6a408f8",
           771 => x"050c82b6",
           772 => x"a408f805",
           773 => x"087082b6",
           774 => x"980c5154",
           775 => x"873d0d82",
           776 => x"b6a40c04",
           777 => x"82b6a408",
           778 => x"0282b6a4",
           779 => x"0ced3d0d",
           780 => x"800b82b6",
           781 => x"a408e405",
           782 => x"2382b6a4",
           783 => x"08880508",
           784 => x"53800b8c",
           785 => x"140c82b6",
           786 => x"a4088805",
           787 => x"08851133",
           788 => x"70812a70",
           789 => x"81327081",
           790 => x"06515151",
           791 => x"51537280",
           792 => x"2e8d38ff",
           793 => x"0b82b6a4",
           794 => x"08e0050c",
           795 => x"96ac3982",
           796 => x"b6a4088c",
           797 => x"05085372",
           798 => x"33537282",
           799 => x"b6a408f8",
           800 => x"05347281",
           801 => x"ff065372",
           802 => x"802e95fa",
           803 => x"3882b6a4",
           804 => x"088c0508",
           805 => x"810582b6",
           806 => x"a4088c05",
           807 => x"0c82b6a4",
           808 => x"08e40522",
           809 => x"70810651",
           810 => x"5372802e",
           811 => x"958b3882",
           812 => x"b6a408f8",
           813 => x"053353af",
           814 => x"732781fc",
           815 => x"3882b6a4",
           816 => x"08f80533",
           817 => x"5372b926",
           818 => x"81ee3882",
           819 => x"b6a408f8",
           820 => x"05335372",
           821 => x"b02e0981",
           822 => x"0680c538",
           823 => x"82b6a408",
           824 => x"e8053370",
           825 => x"982b7098",
           826 => x"2c515153",
           827 => x"72b23882",
           828 => x"b6a408e4",
           829 => x"05227083",
           830 => x"2a708132",
           831 => x"70810651",
           832 => x"51515372",
           833 => x"802e9938",
           834 => x"82b6a408",
           835 => x"e4052270",
           836 => x"82800751",
           837 => x"537282b6",
           838 => x"a408e405",
           839 => x"23fed039",
           840 => x"82b6a408",
           841 => x"e8053370",
           842 => x"982b7098",
           843 => x"2c707083",
           844 => x"2b721173",
           845 => x"11515151",
           846 => x"53515553",
           847 => x"7282b6a4",
           848 => x"08e80534",
           849 => x"82b6a408",
           850 => x"e8053354",
           851 => x"82b6a408",
           852 => x"f8053370",
           853 => x"15d01151",
           854 => x"51537282",
           855 => x"b6a408e8",
           856 => x"053482b6",
           857 => x"a408e805",
           858 => x"3370982b",
           859 => x"70982c51",
           860 => x"51537280",
           861 => x"258b3880",
           862 => x"ff0b82b6",
           863 => x"a408e805",
           864 => x"3482b6a4",
           865 => x"08e40522",
           866 => x"70832a70",
           867 => x"81065151",
           868 => x"5372fddb",
           869 => x"3882b6a4",
           870 => x"08e80533",
           871 => x"70882b70",
           872 => x"902b7090",
           873 => x"2c70882c",
           874 => x"51515151",
           875 => x"537282b6",
           876 => x"a408ec05",
           877 => x"23fdb839",
           878 => x"82b6a408",
           879 => x"e4052270",
           880 => x"832a7081",
           881 => x"06515153",
           882 => x"72802e9d",
           883 => x"3882b6a4",
           884 => x"08e80533",
           885 => x"70982b70",
           886 => x"982c5151",
           887 => x"53728a38",
           888 => x"810b82b6",
           889 => x"a408e805",
           890 => x"3482b6a4",
           891 => x"08f80533",
           892 => x"e01182b6",
           893 => x"a408c405",
           894 => x"0c5382b6",
           895 => x"a408c405",
           896 => x"0880d826",
           897 => x"92943882",
           898 => x"b6a408c4",
           899 => x"05087082",
           900 => x"2b829788",
           901 => x"11700851",
           902 => x"51515372",
           903 => x"0482b6a4",
           904 => x"08e40522",
           905 => x"70900751",
           906 => x"537282b6",
           907 => x"a408e405",
           908 => x"2382b6a4",
           909 => x"08e40522",
           910 => x"70a00751",
           911 => x"537282b6",
           912 => x"a408e405",
           913 => x"23fca839",
           914 => x"82b6a408",
           915 => x"e4052270",
           916 => x"81800751",
           917 => x"537282b6",
           918 => x"a408e405",
           919 => x"23fc9039",
           920 => x"82b6a408",
           921 => x"e4052270",
           922 => x"80c00751",
           923 => x"537282b6",
           924 => x"a408e405",
           925 => x"23fbf839",
           926 => x"82b6a408",
           927 => x"e4052270",
           928 => x"88075153",
           929 => x"7282b6a4",
           930 => x"08e40523",
           931 => x"800b82b6",
           932 => x"a408e805",
           933 => x"34fbd839",
           934 => x"82b6a408",
           935 => x"e4052270",
           936 => x"84075153",
           937 => x"7282b6a4",
           938 => x"08e40523",
           939 => x"fbc139bf",
           940 => x"0b82b6a4",
           941 => x"08fc0534",
           942 => x"82b6a408",
           943 => x"ec0522ff",
           944 => x"11515372",
           945 => x"82b6a408",
           946 => x"ec052380",
           947 => x"e30b82b6",
           948 => x"a408f805",
           949 => x"348da839",
           950 => x"82b6a408",
           951 => x"90050882",
           952 => x"b6a40890",
           953 => x"05088405",
           954 => x"82b6a408",
           955 => x"90050c70",
           956 => x"08515372",
           957 => x"82b6a408",
           958 => x"fc053482",
           959 => x"b6a408ec",
           960 => x"0522ff11",
           961 => x"51537282",
           962 => x"b6a408ec",
           963 => x"05238cef",
           964 => x"3982b6a4",
           965 => x"08900508",
           966 => x"82b6a408",
           967 => x"90050884",
           968 => x"0582b6a4",
           969 => x"0890050c",
           970 => x"700882b6",
           971 => x"a408fc05",
           972 => x"0c82b6a4",
           973 => x"08e40522",
           974 => x"70832a70",
           975 => x"81065151",
           976 => x"51537280",
           977 => x"2eab3882",
           978 => x"b6a408e8",
           979 => x"05337098",
           980 => x"2b537298",
           981 => x"2c5382b6",
           982 => x"a408fc05",
           983 => x"085253a2",
           984 => x"d83f82b6",
           985 => x"98085372",
           986 => x"82b6a408",
           987 => x"f4052399",
           988 => x"3982b6a4",
           989 => x"08fc0508",
           990 => x"519d8a3f",
           991 => x"82b69808",
           992 => x"537282b6",
           993 => x"a408f405",
           994 => x"2382b6a4",
           995 => x"08ec0522",
           996 => x"5382b6a4",
           997 => x"08f40522",
           998 => x"73713154",
           999 => x"547282b6",
          1000 => x"a408ec05",
          1001 => x"238bd839",
          1002 => x"82b6a408",
          1003 => x"90050882",
          1004 => x"b6a40890",
          1005 => x"05088405",
          1006 => x"82b6a408",
          1007 => x"90050c70",
          1008 => x"0882b6a4",
          1009 => x"08fc050c",
          1010 => x"82b6a408",
          1011 => x"e4052270",
          1012 => x"832a7081",
          1013 => x"06515151",
          1014 => x"5372802e",
          1015 => x"ab3882b6",
          1016 => x"a408e805",
          1017 => x"3370982b",
          1018 => x"5372982c",
          1019 => x"5382b6a4",
          1020 => x"08fc0508",
          1021 => x"5253a1c1",
          1022 => x"3f82b698",
          1023 => x"08537282",
          1024 => x"b6a408f4",
          1025 => x"05239939",
          1026 => x"82b6a408",
          1027 => x"fc050851",
          1028 => x"9bf33f82",
          1029 => x"b6980853",
          1030 => x"7282b6a4",
          1031 => x"08f40523",
          1032 => x"82b6a408",
          1033 => x"ec052253",
          1034 => x"82b6a408",
          1035 => x"f4052273",
          1036 => x"71315454",
          1037 => x"7282b6a4",
          1038 => x"08ec0523",
          1039 => x"8ac13982",
          1040 => x"b6a408e4",
          1041 => x"05227082",
          1042 => x"2a708106",
          1043 => x"51515372",
          1044 => x"802ea438",
          1045 => x"82b6a408",
          1046 => x"90050882",
          1047 => x"b6a40890",
          1048 => x"05088405",
          1049 => x"82b6a408",
          1050 => x"90050c70",
          1051 => x"0882b6a4",
          1052 => x"08dc050c",
          1053 => x"53a23982",
          1054 => x"b6a40890",
          1055 => x"050882b6",
          1056 => x"a4089005",
          1057 => x"08840582",
          1058 => x"b6a40890",
          1059 => x"050c7008",
          1060 => x"82b6a408",
          1061 => x"dc050c53",
          1062 => x"82b6a408",
          1063 => x"dc050882",
          1064 => x"b6a408fc",
          1065 => x"050c82b6",
          1066 => x"a408fc05",
          1067 => x"088025a4",
          1068 => x"3882b6a4",
          1069 => x"08e40522",
          1070 => x"70820751",
          1071 => x"537282b6",
          1072 => x"a408e405",
          1073 => x"2382b6a4",
          1074 => x"08fc0508",
          1075 => x"3082b6a4",
          1076 => x"08fc050c",
          1077 => x"82b6a408",
          1078 => x"e4052270",
          1079 => x"ffbf0651",
          1080 => x"537282b6",
          1081 => x"a408e405",
          1082 => x"2381af39",
          1083 => x"880b82b6",
          1084 => x"a408f405",
          1085 => x"23a93982",
          1086 => x"b6a408e4",
          1087 => x"05227080",
          1088 => x"c0075153",
          1089 => x"7282b6a4",
          1090 => x"08e40523",
          1091 => x"80f80b82",
          1092 => x"b6a408f8",
          1093 => x"0534900b",
          1094 => x"82b6a408",
          1095 => x"f4052382",
          1096 => x"b6a408e4",
          1097 => x"05227082",
          1098 => x"2a708106",
          1099 => x"51515372",
          1100 => x"802ea438",
          1101 => x"82b6a408",
          1102 => x"90050882",
          1103 => x"b6a40890",
          1104 => x"05088405",
          1105 => x"82b6a408",
          1106 => x"90050c70",
          1107 => x"0882b6a4",
          1108 => x"08d8050c",
          1109 => x"53a23982",
          1110 => x"b6a40890",
          1111 => x"050882b6",
          1112 => x"a4089005",
          1113 => x"08840582",
          1114 => x"b6a40890",
          1115 => x"050c7008",
          1116 => x"82b6a408",
          1117 => x"d8050c53",
          1118 => x"82b6a408",
          1119 => x"d8050882",
          1120 => x"b6a408fc",
          1121 => x"050c82b6",
          1122 => x"a408e405",
          1123 => x"2270cf06",
          1124 => x"51537282",
          1125 => x"b6a408e4",
          1126 => x"052382b6",
          1127 => x"a80b82b6",
          1128 => x"a408f005",
          1129 => x"0c82b6a4",
          1130 => x"08f00508",
          1131 => x"82b6a408",
          1132 => x"f4052282",
          1133 => x"b6a408fc",
          1134 => x"05087155",
          1135 => x"70545654",
          1136 => x"55a3f33f",
          1137 => x"82b69808",
          1138 => x"53727534",
          1139 => x"82b6a408",
          1140 => x"f0050882",
          1141 => x"b6a408d4",
          1142 => x"050c82b6",
          1143 => x"a408f005",
          1144 => x"08703351",
          1145 => x"53897327",
          1146 => x"a43882b6",
          1147 => x"a408f005",
          1148 => x"08537233",
          1149 => x"5482b6a4",
          1150 => x"08f80533",
          1151 => x"7015df11",
          1152 => x"51515372",
          1153 => x"82b6a408",
          1154 => x"d0053497",
          1155 => x"3982b6a4",
          1156 => x"08f00508",
          1157 => x"537233b0",
          1158 => x"11515372",
          1159 => x"82b6a408",
          1160 => x"d0053482",
          1161 => x"b6a408d4",
          1162 => x"05085382",
          1163 => x"b6a408d0",
          1164 => x"05337334",
          1165 => x"82b6a408",
          1166 => x"f0050881",
          1167 => x"0582b6a4",
          1168 => x"08f0050c",
          1169 => x"82b6a408",
          1170 => x"f4052270",
          1171 => x"5382b6a4",
          1172 => x"08fc0508",
          1173 => x"5253a2ab",
          1174 => x"3f82b698",
          1175 => x"087082b6",
          1176 => x"a408fc05",
          1177 => x"0c5382b6",
          1178 => x"a408fc05",
          1179 => x"08802e84",
          1180 => x"38feb239",
          1181 => x"82b6a408",
          1182 => x"f0050882",
          1183 => x"b6a85455",
          1184 => x"72547470",
          1185 => x"75315153",
          1186 => x"7282b6a4",
          1187 => x"08fc0534",
          1188 => x"82b6a408",
          1189 => x"e4052270",
          1190 => x"b2065153",
          1191 => x"72802e94",
          1192 => x"3882b6a4",
          1193 => x"08ec0522",
          1194 => x"ff115153",
          1195 => x"7282b6a4",
          1196 => x"08ec0523",
          1197 => x"82b6a408",
          1198 => x"e4052270",
          1199 => x"862a7081",
          1200 => x"06515153",
          1201 => x"72802e80",
          1202 => x"e73882b6",
          1203 => x"a408ec05",
          1204 => x"2270902b",
          1205 => x"82b6a408",
          1206 => x"cc050c82",
          1207 => x"b6a408cc",
          1208 => x"0508902c",
          1209 => x"82b6a408",
          1210 => x"cc050c82",
          1211 => x"b6a408f4",
          1212 => x"05225153",
          1213 => x"72902e09",
          1214 => x"81069538",
          1215 => x"82b6a408",
          1216 => x"cc0508fe",
          1217 => x"05537282",
          1218 => x"b6a408c8",
          1219 => x"05239339",
          1220 => x"82b6a408",
          1221 => x"cc0508ff",
          1222 => x"05537282",
          1223 => x"b6a408c8",
          1224 => x"052382b6",
          1225 => x"a408c805",
          1226 => x"2282b6a4",
          1227 => x"08ec0523",
          1228 => x"82b6a408",
          1229 => x"e4052270",
          1230 => x"832a7081",
          1231 => x"06515153",
          1232 => x"72802e80",
          1233 => x"d03882b6",
          1234 => x"a408e805",
          1235 => x"3370982b",
          1236 => x"70982c82",
          1237 => x"b6a408fc",
          1238 => x"05335751",
          1239 => x"51537274",
          1240 => x"24973882",
          1241 => x"b6a408e4",
          1242 => x"052270f7",
          1243 => x"06515372",
          1244 => x"82b6a408",
          1245 => x"e405239d",
          1246 => x"3982b6a4",
          1247 => x"08e80533",
          1248 => x"5382b6a4",
          1249 => x"08fc0533",
          1250 => x"73713154",
          1251 => x"547282b6",
          1252 => x"a408e805",
          1253 => x"3482b6a4",
          1254 => x"08e40522",
          1255 => x"70832a70",
          1256 => x"81065151",
          1257 => x"5372802e",
          1258 => x"b13882b6",
          1259 => x"a408e805",
          1260 => x"3370882b",
          1261 => x"70902b70",
          1262 => x"902c7088",
          1263 => x"2c515151",
          1264 => x"51537254",
          1265 => x"82b6a408",
          1266 => x"ec052270",
          1267 => x"75315153",
          1268 => x"7282b6a4",
          1269 => x"08ec0523",
          1270 => x"af3982b6",
          1271 => x"a408fc05",
          1272 => x"3370882b",
          1273 => x"70902b70",
          1274 => x"902c7088",
          1275 => x"2c515151",
          1276 => x"51537254",
          1277 => x"82b6a408",
          1278 => x"ec052270",
          1279 => x"75315153",
          1280 => x"7282b6a4",
          1281 => x"08ec0523",
          1282 => x"82b6a408",
          1283 => x"e4052270",
          1284 => x"83800651",
          1285 => x"5372b038",
          1286 => x"82b6a408",
          1287 => x"ec0522ff",
          1288 => x"11545472",
          1289 => x"82b6a408",
          1290 => x"ec052373",
          1291 => x"902b7090",
          1292 => x"2c515380",
          1293 => x"73259038",
          1294 => x"82b6a408",
          1295 => x"88050852",
          1296 => x"a0518aee",
          1297 => x"3fd23982",
          1298 => x"b6a408e4",
          1299 => x"05227081",
          1300 => x"2a708106",
          1301 => x"51515372",
          1302 => x"802e9138",
          1303 => x"82b6a408",
          1304 => x"88050852",
          1305 => x"ad518aca",
          1306 => x"3f80c739",
          1307 => x"82b6a408",
          1308 => x"e4052270",
          1309 => x"842a7081",
          1310 => x"06515153",
          1311 => x"72802e90",
          1312 => x"3882b6a4",
          1313 => x"08880508",
          1314 => x"52ab518a",
          1315 => x"a53fa339",
          1316 => x"82b6a408",
          1317 => x"e4052270",
          1318 => x"852a7081",
          1319 => x"06515153",
          1320 => x"72802e8e",
          1321 => x"3882b6a4",
          1322 => x"08880508",
          1323 => x"52a0518a",
          1324 => x"813f82b6",
          1325 => x"a408e405",
          1326 => x"2270862a",
          1327 => x"70810651",
          1328 => x"51537280",
          1329 => x"2eb13882",
          1330 => x"b6a40888",
          1331 => x"050852b0",
          1332 => x"5189df3f",
          1333 => x"82b6a408",
          1334 => x"f4052253",
          1335 => x"72902e09",
          1336 => x"81069438",
          1337 => x"82b6a408",
          1338 => x"88050852",
          1339 => x"82b6a408",
          1340 => x"f8053351",
          1341 => x"89bc3f82",
          1342 => x"b6a408e4",
          1343 => x"05227088",
          1344 => x"2a708106",
          1345 => x"51515372",
          1346 => x"802eb038",
          1347 => x"82b6a408",
          1348 => x"ec0522ff",
          1349 => x"11545472",
          1350 => x"82b6a408",
          1351 => x"ec052373",
          1352 => x"902b7090",
          1353 => x"2c515380",
          1354 => x"73259038",
          1355 => x"82b6a408",
          1356 => x"88050852",
          1357 => x"b05188fa",
          1358 => x"3fd23982",
          1359 => x"b6a408e4",
          1360 => x"05227083",
          1361 => x"2a708106",
          1362 => x"51515372",
          1363 => x"802eb038",
          1364 => x"82b6a408",
          1365 => x"e80533ff",
          1366 => x"11545472",
          1367 => x"82b6a408",
          1368 => x"e8053473",
          1369 => x"982b7098",
          1370 => x"2c515380",
          1371 => x"73259038",
          1372 => x"82b6a408",
          1373 => x"88050852",
          1374 => x"b05188b6",
          1375 => x"3fd23982",
          1376 => x"b6a408e4",
          1377 => x"05227087",
          1378 => x"2a708106",
          1379 => x"51515372",
          1380 => x"b03882b6",
          1381 => x"a408ec05",
          1382 => x"22ff1154",
          1383 => x"547282b6",
          1384 => x"a408ec05",
          1385 => x"2373902b",
          1386 => x"70902c51",
          1387 => x"53807325",
          1388 => x"903882b6",
          1389 => x"a4088805",
          1390 => x"0852a051",
          1391 => x"87f43fd2",
          1392 => x"3982b6a4",
          1393 => x"08f80533",
          1394 => x"537280e3",
          1395 => x"2e098106",
          1396 => x"973882b6",
          1397 => x"a4088805",
          1398 => x"085282b6",
          1399 => x"a408fc05",
          1400 => x"335187ce",
          1401 => x"3f81ee39",
          1402 => x"82b6a408",
          1403 => x"f8053353",
          1404 => x"7280f32e",
          1405 => x"09810680",
          1406 => x"cb3882b6",
          1407 => x"a408f405",
          1408 => x"22ff1151",
          1409 => x"537282b6",
          1410 => x"a408f405",
          1411 => x"237283ff",
          1412 => x"ff065372",
          1413 => x"83ffff2e",
          1414 => x"81bb3882",
          1415 => x"b6a40888",
          1416 => x"05085282",
          1417 => x"b6a408fc",
          1418 => x"05087033",
          1419 => x"5282b6a4",
          1420 => x"08fc0508",
          1421 => x"810582b6",
          1422 => x"a408fc05",
          1423 => x"0c5386f2",
          1424 => x"3fffb739",
          1425 => x"82b6a408",
          1426 => x"f8053353",
          1427 => x"7280d32e",
          1428 => x"09810680",
          1429 => x"cb3882b6",
          1430 => x"a408f405",
          1431 => x"22ff1151",
          1432 => x"537282b6",
          1433 => x"a408f405",
          1434 => x"237283ff",
          1435 => x"ff065372",
          1436 => x"83ffff2e",
          1437 => x"80df3882",
          1438 => x"b6a40888",
          1439 => x"05085282",
          1440 => x"b6a408fc",
          1441 => x"05087033",
          1442 => x"525386a6",
          1443 => x"3f82b6a4",
          1444 => x"08fc0508",
          1445 => x"810582b6",
          1446 => x"a408fc05",
          1447 => x"0cffb739",
          1448 => x"82b6a408",
          1449 => x"f0050882",
          1450 => x"b6a82ea9",
          1451 => x"3882b6a4",
          1452 => x"08880508",
          1453 => x"5282b6a4",
          1454 => x"08f00508",
          1455 => x"ff0582b6",
          1456 => x"a408f005",
          1457 => x"0c82b6a4",
          1458 => x"08f00508",
          1459 => x"70335253",
          1460 => x"85e03fcc",
          1461 => x"3982b6a4",
          1462 => x"08e40522",
          1463 => x"70872a70",
          1464 => x"81065151",
          1465 => x"5372802e",
          1466 => x"80c33882",
          1467 => x"b6a408ec",
          1468 => x"0522ff11",
          1469 => x"54547282",
          1470 => x"b6a408ec",
          1471 => x"05237390",
          1472 => x"2b70902c",
          1473 => x"51538073",
          1474 => x"25a33882",
          1475 => x"b6a40888",
          1476 => x"050852a0",
          1477 => x"51859b3f",
          1478 => x"d23982b6",
          1479 => x"a4088805",
          1480 => x"085282b6",
          1481 => x"a408f805",
          1482 => x"33518586",
          1483 => x"3f800b82",
          1484 => x"b6a408e4",
          1485 => x"0523eab7",
          1486 => x"3982b6a4",
          1487 => x"08f80533",
          1488 => x"5372a52e",
          1489 => x"098106a8",
          1490 => x"38810b82",
          1491 => x"b6a408e4",
          1492 => x"0523800b",
          1493 => x"82b6a408",
          1494 => x"ec052380",
          1495 => x"0b82b6a4",
          1496 => x"08e80534",
          1497 => x"8a0b82b6",
          1498 => x"a408f405",
          1499 => x"23ea8039",
          1500 => x"82b6a408",
          1501 => x"88050852",
          1502 => x"82b6a408",
          1503 => x"f8053351",
          1504 => x"84b03fe9",
          1505 => x"ea3982b6",
          1506 => x"a4088805",
          1507 => x"088c1108",
          1508 => x"7082b6a4",
          1509 => x"08e0050c",
          1510 => x"515382b6",
          1511 => x"a408e005",
          1512 => x"0882b698",
          1513 => x"0c953d0d",
          1514 => x"82b6a40c",
          1515 => x"0482b6a4",
          1516 => x"080282b6",
          1517 => x"a40cfd3d",
          1518 => x"0d82cde8",
          1519 => x"085382b6",
          1520 => x"a4088c05",
          1521 => x"085282b6",
          1522 => x"a4088805",
          1523 => x"0851e4dd",
          1524 => x"3f82b698",
          1525 => x"087082b6",
          1526 => x"980c5485",
          1527 => x"3d0d82b6",
          1528 => x"a40c0482",
          1529 => x"b6a40802",
          1530 => x"82b6a40c",
          1531 => x"fb3d0d80",
          1532 => x"0b82b6a4",
          1533 => x"08f8050c",
          1534 => x"82cdec08",
          1535 => x"85113370",
          1536 => x"812a7081",
          1537 => x"32708106",
          1538 => x"51515151",
          1539 => x"5372802e",
          1540 => x"8d38ff0b",
          1541 => x"82b6a408",
          1542 => x"f4050c81",
          1543 => x"923982b6",
          1544 => x"a4088805",
          1545 => x"08537233",
          1546 => x"82b6a408",
          1547 => x"88050881",
          1548 => x"0582b6a4",
          1549 => x"0888050c",
          1550 => x"537282b6",
          1551 => x"a408fc05",
          1552 => x"347281ff",
          1553 => x"06537280",
          1554 => x"2eb03882",
          1555 => x"cdec0882",
          1556 => x"cdec0853",
          1557 => x"82b6a408",
          1558 => x"fc053352",
          1559 => x"90110851",
          1560 => x"53722d82",
          1561 => x"b6980853",
          1562 => x"72802eff",
          1563 => x"b138ff0b",
          1564 => x"82b6a408",
          1565 => x"f8050cff",
          1566 => x"a53982cd",
          1567 => x"ec0882cd",
          1568 => x"ec085353",
          1569 => x"8a519013",
          1570 => x"0853722d",
          1571 => x"82b69808",
          1572 => x"5372802e",
          1573 => x"8a38ff0b",
          1574 => x"82b6a408",
          1575 => x"f8050c82",
          1576 => x"b6a408f8",
          1577 => x"05087082",
          1578 => x"b6a408f4",
          1579 => x"050c5382",
          1580 => x"b6a408f4",
          1581 => x"050882b6",
          1582 => x"980c873d",
          1583 => x"0d82b6a4",
          1584 => x"0c0482b6",
          1585 => x"a4080282",
          1586 => x"b6a40cfb",
          1587 => x"3d0d800b",
          1588 => x"82b6a408",
          1589 => x"f8050c82",
          1590 => x"b6a4088c",
          1591 => x"05088511",
          1592 => x"3370812a",
          1593 => x"70813270",
          1594 => x"81065151",
          1595 => x"51515372",
          1596 => x"802e8d38",
          1597 => x"ff0b82b6",
          1598 => x"a408f405",
          1599 => x"0c80f339",
          1600 => x"82b6a408",
          1601 => x"88050853",
          1602 => x"723382b6",
          1603 => x"a4088805",
          1604 => x"08810582",
          1605 => x"b6a40888",
          1606 => x"050c5372",
          1607 => x"82b6a408",
          1608 => x"fc053472",
          1609 => x"81ff0653",
          1610 => x"72802eb6",
          1611 => x"3882b6a4",
          1612 => x"088c0508",
          1613 => x"82b6a408",
          1614 => x"8c050853",
          1615 => x"82b6a408",
          1616 => x"fc053352",
          1617 => x"90110851",
          1618 => x"53722d82",
          1619 => x"b6980853",
          1620 => x"72802eff",
          1621 => x"ab38ff0b",
          1622 => x"82b6a408",
          1623 => x"f8050cff",
          1624 => x"9f3982b6",
          1625 => x"a408f805",
          1626 => x"087082b6",
          1627 => x"a408f405",
          1628 => x"0c5382b6",
          1629 => x"a408f405",
          1630 => x"0882b698",
          1631 => x"0c873d0d",
          1632 => x"82b6a40c",
          1633 => x"0482b6a4",
          1634 => x"080282b6",
          1635 => x"a40cfe3d",
          1636 => x"0d82cdec",
          1637 => x"085282b6",
          1638 => x"a4088805",
          1639 => x"0851933f",
          1640 => x"82b69808",
          1641 => x"7082b698",
          1642 => x"0c53843d",
          1643 => x"0d82b6a4",
          1644 => x"0c0482b6",
          1645 => x"a4080282",
          1646 => x"b6a40cfb",
          1647 => x"3d0d82b6",
          1648 => x"a4088c05",
          1649 => x"08851133",
          1650 => x"70812a70",
          1651 => x"81327081",
          1652 => x"06515151",
          1653 => x"51537280",
          1654 => x"2e8d38ff",
          1655 => x"0b82b6a4",
          1656 => x"08fc050c",
          1657 => x"81cb3982",
          1658 => x"b6a4088c",
          1659 => x"05088511",
          1660 => x"3370822a",
          1661 => x"70810651",
          1662 => x"51515372",
          1663 => x"802e80db",
          1664 => x"3882b6a4",
          1665 => x"088c0508",
          1666 => x"82b6a408",
          1667 => x"8c050854",
          1668 => x"548c1408",
          1669 => x"88140825",
          1670 => x"9f3882b6",
          1671 => x"a4088c05",
          1672 => x"08700870",
          1673 => x"82b6a408",
          1674 => x"88050852",
          1675 => x"57545472",
          1676 => x"75347308",
          1677 => x"8105740c",
          1678 => x"82b6a408",
          1679 => x"8c05088c",
          1680 => x"11088105",
          1681 => x"8c120c82",
          1682 => x"b6a40888",
          1683 => x"05087082",
          1684 => x"b6a408fc",
          1685 => x"050c5153",
          1686 => x"80d73982",
          1687 => x"b6a4088c",
          1688 => x"050882b6",
          1689 => x"a4088c05",
          1690 => x"085382b6",
          1691 => x"a4088805",
          1692 => x"087081ff",
          1693 => x"06539012",
          1694 => x"08515454",
          1695 => x"722d82b6",
          1696 => x"98085372",
          1697 => x"a33882b6",
          1698 => x"a4088c05",
          1699 => x"088c1108",
          1700 => x"81058c12",
          1701 => x"0c82b6a4",
          1702 => x"08880508",
          1703 => x"7082b6a4",
          1704 => x"08fc050c",
          1705 => x"51538a39",
          1706 => x"ff0b82b6",
          1707 => x"a408fc05",
          1708 => x"0c82b6a4",
          1709 => x"08fc0508",
          1710 => x"82b6980c",
          1711 => x"873d0d82",
          1712 => x"b6a40c04",
          1713 => x"82b6a408",
          1714 => x"0282b6a4",
          1715 => x"0cf93d0d",
          1716 => x"82b6a408",
          1717 => x"88050885",
          1718 => x"11337081",
          1719 => x"32708106",
          1720 => x"51515152",
          1721 => x"71802e8d",
          1722 => x"38ff0b82",
          1723 => x"b6a408f8",
          1724 => x"050c8394",
          1725 => x"3982b6a4",
          1726 => x"08880508",
          1727 => x"85113370",
          1728 => x"862a7081",
          1729 => x"06515151",
          1730 => x"5271802e",
          1731 => x"80c53882",
          1732 => x"b6a40888",
          1733 => x"050882b6",
          1734 => x"a4088805",
          1735 => x"08535385",
          1736 => x"123370ff",
          1737 => x"bf065152",
          1738 => x"71851434",
          1739 => x"82b6a408",
          1740 => x"8805088c",
          1741 => x"11088105",
          1742 => x"8c120c82",
          1743 => x"b6a40888",
          1744 => x"05088411",
          1745 => x"337082b6",
          1746 => x"a408f805",
          1747 => x"0c515152",
          1748 => x"82b63982",
          1749 => x"b6a40888",
          1750 => x"05088511",
          1751 => x"3370822a",
          1752 => x"70810651",
          1753 => x"51515271",
          1754 => x"802e80d7",
          1755 => x"3882b6a4",
          1756 => x"08880508",
          1757 => x"70087033",
          1758 => x"82b6a408",
          1759 => x"fc050c51",
          1760 => x"5282b6a4",
          1761 => x"08fc0508",
          1762 => x"a93882b6",
          1763 => x"a4088805",
          1764 => x"0882b6a4",
          1765 => x"08880508",
          1766 => x"53538512",
          1767 => x"3370a007",
          1768 => x"51527185",
          1769 => x"1434ff0b",
          1770 => x"82b6a408",
          1771 => x"f8050c81",
          1772 => x"d73982b6",
          1773 => x"a4088805",
          1774 => x"08700881",
          1775 => x"05710c52",
          1776 => x"81a13982",
          1777 => x"b6a40888",
          1778 => x"050882b6",
          1779 => x"a4088805",
          1780 => x"08529411",
          1781 => x"08515271",
          1782 => x"2d82b698",
          1783 => x"087082b6",
          1784 => x"a408fc05",
          1785 => x"0c5282b6",
          1786 => x"a408fc05",
          1787 => x"08802580",
          1788 => x"f23882b6",
          1789 => x"a4088805",
          1790 => x"0882b6a4",
          1791 => x"08f4050c",
          1792 => x"82b6a408",
          1793 => x"88050885",
          1794 => x"113382b6",
          1795 => x"a408f005",
          1796 => x"0c5282b6",
          1797 => x"a408fc05",
          1798 => x"08ff2e09",
          1799 => x"81069538",
          1800 => x"82b6a408",
          1801 => x"f0050890",
          1802 => x"07527182",
          1803 => x"b6a408ec",
          1804 => x"05349339",
          1805 => x"82b6a408",
          1806 => x"f00508a0",
          1807 => x"07527182",
          1808 => x"b6a408ec",
          1809 => x"053482b6",
          1810 => x"a408f405",
          1811 => x"085282b6",
          1812 => x"a408ec05",
          1813 => x"33851334",
          1814 => x"ff0b82b6",
          1815 => x"a408f805",
          1816 => x"0ca63982",
          1817 => x"b6a40888",
          1818 => x"05088c11",
          1819 => x"0881058c",
          1820 => x"120c82b6",
          1821 => x"a408fc05",
          1822 => x"087081ff",
          1823 => x"067082b6",
          1824 => x"a408f805",
          1825 => x"0c515152",
          1826 => x"82b6a408",
          1827 => x"f8050882",
          1828 => x"b6980c89",
          1829 => x"3d0d82b6",
          1830 => x"a40c0482",
          1831 => x"b6a40802",
          1832 => x"82b6a40c",
          1833 => x"fd3d0d82",
          1834 => x"b6a40888",
          1835 => x"050882b6",
          1836 => x"a408fc05",
          1837 => x"0c82b6a4",
          1838 => x"088c0508",
          1839 => x"82b6a408",
          1840 => x"f8050c82",
          1841 => x"b6a40890",
          1842 => x"0508802e",
          1843 => x"82a23882",
          1844 => x"b6a408f8",
          1845 => x"050882b6",
          1846 => x"a408fc05",
          1847 => x"082681ac",
          1848 => x"3882b6a4",
          1849 => x"08f80508",
          1850 => x"82b6a408",
          1851 => x"90050805",
          1852 => x"5182b6a4",
          1853 => x"08fc0508",
          1854 => x"71278190",
          1855 => x"3882b6a4",
          1856 => x"08fc0508",
          1857 => x"82b6a408",
          1858 => x"90050805",
          1859 => x"82b6a408",
          1860 => x"fc050c82",
          1861 => x"b6a408f8",
          1862 => x"050882b6",
          1863 => x"a4089005",
          1864 => x"080582b6",
          1865 => x"a408f805",
          1866 => x"0c82b6a4",
          1867 => x"08900508",
          1868 => x"810582b6",
          1869 => x"a4089005",
          1870 => x"0c82b6a4",
          1871 => x"08900508",
          1872 => x"ff0582b6",
          1873 => x"a4089005",
          1874 => x"0c82b6a4",
          1875 => x"08900508",
          1876 => x"802e819c",
          1877 => x"3882b6a4",
          1878 => x"08fc0508",
          1879 => x"ff0582b6",
          1880 => x"a408fc05",
          1881 => x"0c82b6a4",
          1882 => x"08f80508",
          1883 => x"ff0582b6",
          1884 => x"a408f805",
          1885 => x"0c82b6a4",
          1886 => x"08fc0508",
          1887 => x"82b6a408",
          1888 => x"f8050853",
          1889 => x"51713371",
          1890 => x"34ffae39",
          1891 => x"82b6a408",
          1892 => x"90050881",
          1893 => x"0582b6a4",
          1894 => x"0890050c",
          1895 => x"82b6a408",
          1896 => x"900508ff",
          1897 => x"0582b6a4",
          1898 => x"0890050c",
          1899 => x"82b6a408",
          1900 => x"90050880",
          1901 => x"2eba3882",
          1902 => x"b6a408f8",
          1903 => x"05085170",
          1904 => x"3382b6a4",
          1905 => x"08f80508",
          1906 => x"810582b6",
          1907 => x"a408f805",
          1908 => x"0c82b6a4",
          1909 => x"08fc0508",
          1910 => x"52527171",
          1911 => x"3482b6a4",
          1912 => x"08fc0508",
          1913 => x"810582b6",
          1914 => x"a408fc05",
          1915 => x"0cffad39",
          1916 => x"82b6a408",
          1917 => x"88050870",
          1918 => x"82b6980c",
          1919 => x"51853d0d",
          1920 => x"82b6a40c",
          1921 => x"0482b6a4",
          1922 => x"080282b6",
          1923 => x"a40cfe3d",
          1924 => x"0d82b6a4",
          1925 => x"08880508",
          1926 => x"82b6a408",
          1927 => x"fc050c82",
          1928 => x"b6a408fc",
          1929 => x"05085271",
          1930 => x"3382b6a4",
          1931 => x"08fc0508",
          1932 => x"810582b6",
          1933 => x"a408fc05",
          1934 => x"0c7081ff",
          1935 => x"06515170",
          1936 => x"802e8338",
          1937 => x"da3982b6",
          1938 => x"a408fc05",
          1939 => x"08ff0582",
          1940 => x"b6a408fc",
          1941 => x"050c82b6",
          1942 => x"a408fc05",
          1943 => x"0882b6a4",
          1944 => x"08880508",
          1945 => x"317082b6",
          1946 => x"980c5184",
          1947 => x"3d0d82b6",
          1948 => x"a40c0482",
          1949 => x"b6a40802",
          1950 => x"82b6a40c",
          1951 => x"fe3d0d82",
          1952 => x"b6a40888",
          1953 => x"050882b6",
          1954 => x"a408fc05",
          1955 => x"0c82b6a4",
          1956 => x"088c0508",
          1957 => x"52713382",
          1958 => x"b6a4088c",
          1959 => x"05088105",
          1960 => x"82b6a408",
          1961 => x"8c050c82",
          1962 => x"b6a408fc",
          1963 => x"05085351",
          1964 => x"70723482",
          1965 => x"b6a408fc",
          1966 => x"05088105",
          1967 => x"82b6a408",
          1968 => x"fc050c70",
          1969 => x"81ff0651",
          1970 => x"70802e84",
          1971 => x"38ffbe39",
          1972 => x"82b6a408",
          1973 => x"88050870",
          1974 => x"82b6980c",
          1975 => x"51843d0d",
          1976 => x"82b6a40c",
          1977 => x"0482b6a4",
          1978 => x"080282b6",
          1979 => x"a40cfd3d",
          1980 => x"0d82b6a4",
          1981 => x"08880508",
          1982 => x"82b6a408",
          1983 => x"fc050c82",
          1984 => x"b6a4088c",
          1985 => x"050882b6",
          1986 => x"a408f805",
          1987 => x"0c82b6a4",
          1988 => x"08900508",
          1989 => x"802e80e5",
          1990 => x"3882b6a4",
          1991 => x"08900508",
          1992 => x"810582b6",
          1993 => x"a4089005",
          1994 => x"0c82b6a4",
          1995 => x"08900508",
          1996 => x"ff0582b6",
          1997 => x"a4089005",
          1998 => x"0c82b6a4",
          1999 => x"08900508",
          2000 => x"802eba38",
          2001 => x"82b6a408",
          2002 => x"f8050851",
          2003 => x"703382b6",
          2004 => x"a408f805",
          2005 => x"08810582",
          2006 => x"b6a408f8",
          2007 => x"050c82b6",
          2008 => x"a408fc05",
          2009 => x"08525271",
          2010 => x"713482b6",
          2011 => x"a408fc05",
          2012 => x"08810582",
          2013 => x"b6a408fc",
          2014 => x"050cffad",
          2015 => x"3982b6a4",
          2016 => x"08880508",
          2017 => x"7082b698",
          2018 => x"0c51853d",
          2019 => x"0d82b6a4",
          2020 => x"0c0482b6",
          2021 => x"a4080282",
          2022 => x"b6a40cfd",
          2023 => x"3d0d82b6",
          2024 => x"a4089005",
          2025 => x"08802e81",
          2026 => x"f43882b6",
          2027 => x"a4088c05",
          2028 => x"08527133",
          2029 => x"82b6a408",
          2030 => x"8c050881",
          2031 => x"0582b6a4",
          2032 => x"088c050c",
          2033 => x"82b6a408",
          2034 => x"88050870",
          2035 => x"337281ff",
          2036 => x"06535454",
          2037 => x"5171712e",
          2038 => x"843880ce",
          2039 => x"3982b6a4",
          2040 => x"08880508",
          2041 => x"52713382",
          2042 => x"b6a40888",
          2043 => x"05088105",
          2044 => x"82b6a408",
          2045 => x"88050c70",
          2046 => x"81ff0651",
          2047 => x"51708d38",
          2048 => x"800b82b6",
          2049 => x"a408fc05",
          2050 => x"0c819b39",
          2051 => x"82b6a408",
          2052 => x"900508ff",
          2053 => x"0582b6a4",
          2054 => x"0890050c",
          2055 => x"82b6a408",
          2056 => x"90050880",
          2057 => x"2e8438ff",
          2058 => x"813982b6",
          2059 => x"a4089005",
          2060 => x"08802e80",
          2061 => x"e83882b6",
          2062 => x"a4088805",
          2063 => x"08703352",
          2064 => x"53708d38",
          2065 => x"ff0b82b6",
          2066 => x"a408fc05",
          2067 => x"0c80d739",
          2068 => x"82b6a408",
          2069 => x"8c0508ff",
          2070 => x"0582b6a4",
          2071 => x"088c050c",
          2072 => x"82b6a408",
          2073 => x"8c050870",
          2074 => x"33525270",
          2075 => x"8c38810b",
          2076 => x"82b6a408",
          2077 => x"fc050cae",
          2078 => x"3982b6a4",
          2079 => x"08880508",
          2080 => x"703382b6",
          2081 => x"a4088c05",
          2082 => x"08703372",
          2083 => x"71317082",
          2084 => x"b6a408fc",
          2085 => x"050c5355",
          2086 => x"5252538a",
          2087 => x"39800b82",
          2088 => x"b6a408fc",
          2089 => x"050c82b6",
          2090 => x"a408fc05",
          2091 => x"0882b698",
          2092 => x"0c853d0d",
          2093 => x"82b6a40c",
          2094 => x"0482b6a4",
          2095 => x"080282b6",
          2096 => x"a40cfd3d",
          2097 => x"0d82b6a4",
          2098 => x"08880508",
          2099 => x"82b6a408",
          2100 => x"f8050c82",
          2101 => x"b6a4088c",
          2102 => x"05088d38",
          2103 => x"800b82b6",
          2104 => x"a408fc05",
          2105 => x"0c80ec39",
          2106 => x"82b6a408",
          2107 => x"f8050852",
          2108 => x"713382b6",
          2109 => x"a408f805",
          2110 => x"08810582",
          2111 => x"b6a408f8",
          2112 => x"050c7081",
          2113 => x"ff065151",
          2114 => x"70802e9f",
          2115 => x"3882b6a4",
          2116 => x"088c0508",
          2117 => x"ff0582b6",
          2118 => x"a4088c05",
          2119 => x"0c82b6a4",
          2120 => x"088c0508",
          2121 => x"ff2e8438",
          2122 => x"ffbe3982",
          2123 => x"b6a408f8",
          2124 => x"0508ff05",
          2125 => x"82b6a408",
          2126 => x"f8050c82",
          2127 => x"b6a408f8",
          2128 => x"050882b6",
          2129 => x"a4088805",
          2130 => x"08317082",
          2131 => x"b6a408fc",
          2132 => x"050c5182",
          2133 => x"b6a408fc",
          2134 => x"050882b6",
          2135 => x"980c853d",
          2136 => x"0d82b6a4",
          2137 => x"0c0482b6",
          2138 => x"a4080282",
          2139 => x"b6a40cfe",
          2140 => x"3d0d82b6",
          2141 => x"a4088805",
          2142 => x"0882b6a4",
          2143 => x"08fc050c",
          2144 => x"82b6a408",
          2145 => x"90050880",
          2146 => x"2e80d438",
          2147 => x"82b6a408",
          2148 => x"90050881",
          2149 => x"0582b6a4",
          2150 => x"0890050c",
          2151 => x"82b6a408",
          2152 => x"900508ff",
          2153 => x"0582b6a4",
          2154 => x"0890050c",
          2155 => x"82b6a408",
          2156 => x"90050880",
          2157 => x"2ea93882",
          2158 => x"b6a4088c",
          2159 => x"05085170",
          2160 => x"82b6a408",
          2161 => x"fc050852",
          2162 => x"52717134",
          2163 => x"82b6a408",
          2164 => x"fc050881",
          2165 => x"0582b6a4",
          2166 => x"08fc050c",
          2167 => x"ffbe3982",
          2168 => x"b6a40888",
          2169 => x"05087082",
          2170 => x"b6980c51",
          2171 => x"843d0d82",
          2172 => x"b6a40c04",
          2173 => x"82b6a408",
          2174 => x"0282b6a4",
          2175 => x"0cf93d0d",
          2176 => x"800b82b6",
          2177 => x"a408fc05",
          2178 => x"0c82b6a4",
          2179 => x"08880508",
          2180 => x"8025b938",
          2181 => x"82b6a408",
          2182 => x"88050830",
          2183 => x"82b6a408",
          2184 => x"88050c80",
          2185 => x"0b82b6a4",
          2186 => x"08f4050c",
          2187 => x"82b6a408",
          2188 => x"fc05088a",
          2189 => x"38810b82",
          2190 => x"b6a408f4",
          2191 => x"050c82b6",
          2192 => x"a408f405",
          2193 => x"0882b6a4",
          2194 => x"08fc050c",
          2195 => x"82b6a408",
          2196 => x"8c050880",
          2197 => x"25b93882",
          2198 => x"b6a4088c",
          2199 => x"05083082",
          2200 => x"b6a4088c",
          2201 => x"050c800b",
          2202 => x"82b6a408",
          2203 => x"f0050c82",
          2204 => x"b6a408fc",
          2205 => x"05088a38",
          2206 => x"810b82b6",
          2207 => x"a408f005",
          2208 => x"0c82b6a4",
          2209 => x"08f00508",
          2210 => x"82b6a408",
          2211 => x"fc050c80",
          2212 => x"5382b6a4",
          2213 => x"088c0508",
          2214 => x"5282b6a4",
          2215 => x"08880508",
          2216 => x"5182c53f",
          2217 => x"82b69808",
          2218 => x"7082b6a4",
          2219 => x"08f8050c",
          2220 => x"5482b6a4",
          2221 => x"08fc0508",
          2222 => x"802e9038",
          2223 => x"82b6a408",
          2224 => x"f8050830",
          2225 => x"82b6a408",
          2226 => x"f8050c82",
          2227 => x"b6a408f8",
          2228 => x"05087082",
          2229 => x"b6980c54",
          2230 => x"893d0d82",
          2231 => x"b6a40c04",
          2232 => x"82b6a408",
          2233 => x"0282b6a4",
          2234 => x"0cfb3d0d",
          2235 => x"800b82b6",
          2236 => x"a408fc05",
          2237 => x"0c82b6a4",
          2238 => x"08880508",
          2239 => x"80259938",
          2240 => x"82b6a408",
          2241 => x"88050830",
          2242 => x"82b6a408",
          2243 => x"88050c81",
          2244 => x"0b82b6a4",
          2245 => x"08fc050c",
          2246 => x"82b6a408",
          2247 => x"8c050880",
          2248 => x"25903882",
          2249 => x"b6a4088c",
          2250 => x"05083082",
          2251 => x"b6a4088c",
          2252 => x"050c8153",
          2253 => x"82b6a408",
          2254 => x"8c050852",
          2255 => x"82b6a408",
          2256 => x"88050851",
          2257 => x"81a23f82",
          2258 => x"b6980870",
          2259 => x"82b6a408",
          2260 => x"f8050c54",
          2261 => x"82b6a408",
          2262 => x"fc050880",
          2263 => x"2e903882",
          2264 => x"b6a408f8",
          2265 => x"05083082",
          2266 => x"b6a408f8",
          2267 => x"050c82b6",
          2268 => x"a408f805",
          2269 => x"087082b6",
          2270 => x"980c5487",
          2271 => x"3d0d82b6",
          2272 => x"a40c0482",
          2273 => x"b6a40802",
          2274 => x"82b6a40c",
          2275 => x"fd3d0d80",
          2276 => x"5382b6a4",
          2277 => x"088c0508",
          2278 => x"5282b6a4",
          2279 => x"08880508",
          2280 => x"5180c53f",
          2281 => x"82b69808",
          2282 => x"7082b698",
          2283 => x"0c54853d",
          2284 => x"0d82b6a4",
          2285 => x"0c0482b6",
          2286 => x"a4080282",
          2287 => x"b6a40cfd",
          2288 => x"3d0d8153",
          2289 => x"82b6a408",
          2290 => x"8c050852",
          2291 => x"82b6a408",
          2292 => x"88050851",
          2293 => x"933f82b6",
          2294 => x"98087082",
          2295 => x"b6980c54",
          2296 => x"853d0d82",
          2297 => x"b6a40c04",
          2298 => x"82b6a408",
          2299 => x"0282b6a4",
          2300 => x"0cfd3d0d",
          2301 => x"810b82b6",
          2302 => x"a408fc05",
          2303 => x"0c800b82",
          2304 => x"b6a408f8",
          2305 => x"050c82b6",
          2306 => x"a4088c05",
          2307 => x"0882b6a4",
          2308 => x"08880508",
          2309 => x"27b93882",
          2310 => x"b6a408fc",
          2311 => x"0508802e",
          2312 => x"ae38800b",
          2313 => x"82b6a408",
          2314 => x"8c050824",
          2315 => x"a23882b6",
          2316 => x"a4088c05",
          2317 => x"081082b6",
          2318 => x"a4088c05",
          2319 => x"0c82b6a4",
          2320 => x"08fc0508",
          2321 => x"1082b6a4",
          2322 => x"08fc050c",
          2323 => x"ffb83982",
          2324 => x"b6a408fc",
          2325 => x"0508802e",
          2326 => x"80e13882",
          2327 => x"b6a4088c",
          2328 => x"050882b6",
          2329 => x"a4088805",
          2330 => x"0826ad38",
          2331 => x"82b6a408",
          2332 => x"88050882",
          2333 => x"b6a4088c",
          2334 => x"05083182",
          2335 => x"b6a40888",
          2336 => x"050c82b6",
          2337 => x"a408f805",
          2338 => x"0882b6a4",
          2339 => x"08fc0508",
          2340 => x"0782b6a4",
          2341 => x"08f8050c",
          2342 => x"82b6a408",
          2343 => x"fc050881",
          2344 => x"2a82b6a4",
          2345 => x"08fc050c",
          2346 => x"82b6a408",
          2347 => x"8c050881",
          2348 => x"2a82b6a4",
          2349 => x"088c050c",
          2350 => x"ff953982",
          2351 => x"b6a40890",
          2352 => x"0508802e",
          2353 => x"933882b6",
          2354 => x"a4088805",
          2355 => x"087082b6",
          2356 => x"a408f405",
          2357 => x"0c519139",
          2358 => x"82b6a408",
          2359 => x"f8050870",
          2360 => x"82b6a408",
          2361 => x"f4050c51",
          2362 => x"82b6a408",
          2363 => x"f4050882",
          2364 => x"b6980c85",
          2365 => x"3d0d82b6",
          2366 => x"a40c0482",
          2367 => x"b6a40802",
          2368 => x"82b6a40c",
          2369 => x"f73d0d80",
          2370 => x"0b82b6a4",
          2371 => x"08f00534",
          2372 => x"82b6a408",
          2373 => x"8c050853",
          2374 => x"80730c82",
          2375 => x"b6a40888",
          2376 => x"05087008",
          2377 => x"51537233",
          2378 => x"537282b6",
          2379 => x"a408f805",
          2380 => x"347281ff",
          2381 => x"065372a0",
          2382 => x"2e098106",
          2383 => x"913882b6",
          2384 => x"a4088805",
          2385 => x"08700881",
          2386 => x"05710c53",
          2387 => x"ce3982b6",
          2388 => x"a408f805",
          2389 => x"335372ad",
          2390 => x"2e098106",
          2391 => x"a438810b",
          2392 => x"82b6a408",
          2393 => x"f0053482",
          2394 => x"b6a40888",
          2395 => x"05087008",
          2396 => x"8105710c",
          2397 => x"70085153",
          2398 => x"723382b6",
          2399 => x"a408f805",
          2400 => x"3482b6a4",
          2401 => x"08f80533",
          2402 => x"5372b02e",
          2403 => x"09810681",
          2404 => x"dc3882b6",
          2405 => x"a4088805",
          2406 => x"08700881",
          2407 => x"05710c70",
          2408 => x"08515372",
          2409 => x"3382b6a4",
          2410 => x"08f80534",
          2411 => x"82b6a408",
          2412 => x"f8053382",
          2413 => x"b6a408e8",
          2414 => x"050c82b6",
          2415 => x"a408e805",
          2416 => x"0880e22e",
          2417 => x"b63882b6",
          2418 => x"a408e805",
          2419 => x"0880f82e",
          2420 => x"843880cd",
          2421 => x"39900b82",
          2422 => x"b6a408f4",
          2423 => x"053482b6",
          2424 => x"a4088805",
          2425 => x"08700881",
          2426 => x"05710c70",
          2427 => x"08515372",
          2428 => x"3382b6a4",
          2429 => x"08f80534",
          2430 => x"81a43982",
          2431 => x"0b82b6a4",
          2432 => x"08f40534",
          2433 => x"82b6a408",
          2434 => x"88050870",
          2435 => x"08810571",
          2436 => x"0c700851",
          2437 => x"53723382",
          2438 => x"b6a408f8",
          2439 => x"053480fe",
          2440 => x"3982b6a4",
          2441 => x"08f80533",
          2442 => x"5372a026",
          2443 => x"8d38810b",
          2444 => x"82b6a408",
          2445 => x"ec050c83",
          2446 => x"803982b6",
          2447 => x"a408f805",
          2448 => x"3353af73",
          2449 => x"27903882",
          2450 => x"b6a408f8",
          2451 => x"05335372",
          2452 => x"b9268338",
          2453 => x"8d39800b",
          2454 => x"82b6a408",
          2455 => x"ec050c82",
          2456 => x"d839880b",
          2457 => x"82b6a408",
          2458 => x"f40534b2",
          2459 => x"3982b6a4",
          2460 => x"08f80533",
          2461 => x"53af7327",
          2462 => x"903882b6",
          2463 => x"a408f805",
          2464 => x"335372b9",
          2465 => x"2683388d",
          2466 => x"39800b82",
          2467 => x"b6a408ec",
          2468 => x"050c82a5",
          2469 => x"398a0b82",
          2470 => x"b6a408f4",
          2471 => x"0534800b",
          2472 => x"82b6a408",
          2473 => x"fc050c82",
          2474 => x"b6a408f8",
          2475 => x"053353a0",
          2476 => x"732781cf",
          2477 => x"3882b6a4",
          2478 => x"08f80533",
          2479 => x"5380e073",
          2480 => x"27943882",
          2481 => x"b6a408f8",
          2482 => x"0533e011",
          2483 => x"51537282",
          2484 => x"b6a408f8",
          2485 => x"053482b6",
          2486 => x"a408f805",
          2487 => x"33d01151",
          2488 => x"537282b6",
          2489 => x"a408f805",
          2490 => x"3482b6a4",
          2491 => x"08f80533",
          2492 => x"53907327",
          2493 => x"ad3882b6",
          2494 => x"a408f805",
          2495 => x"33f91151",
          2496 => x"537282b6",
          2497 => x"a408f805",
          2498 => x"3482b6a4",
          2499 => x"08f80533",
          2500 => x"53728926",
          2501 => x"8d38800b",
          2502 => x"82b6a408",
          2503 => x"ec050c81",
          2504 => x"983982b6",
          2505 => x"a408f805",
          2506 => x"3382b6a4",
          2507 => x"08f40533",
          2508 => x"54547274",
          2509 => x"268d3880",
          2510 => x"0b82b6a4",
          2511 => x"08ec050c",
          2512 => x"80f73982",
          2513 => x"b6a408f4",
          2514 => x"05337082",
          2515 => x"b6a408fc",
          2516 => x"05082982",
          2517 => x"b6a408f8",
          2518 => x"05337012",
          2519 => x"82b6a408",
          2520 => x"fc050c82",
          2521 => x"b6a40888",
          2522 => x"05087008",
          2523 => x"8105710c",
          2524 => x"70085151",
          2525 => x"52555372",
          2526 => x"3382b6a4",
          2527 => x"08f80534",
          2528 => x"fea53982",
          2529 => x"b6a408f0",
          2530 => x"05335372",
          2531 => x"802e9038",
          2532 => x"82b6a408",
          2533 => x"fc050830",
          2534 => x"82b6a408",
          2535 => x"fc050c82",
          2536 => x"b6a4088c",
          2537 => x"050882b6",
          2538 => x"a408fc05",
          2539 => x"08710c53",
          2540 => x"810b82b6",
          2541 => x"a408ec05",
          2542 => x"0c82b6a4",
          2543 => x"08ec0508",
          2544 => x"82b6980c",
          2545 => x"8b3d0d82",
          2546 => x"b6a40c04",
          2547 => x"82b6a408",
          2548 => x"0282b6a4",
          2549 => x"0cf73d0d",
          2550 => x"800b82b6",
          2551 => x"a408f005",
          2552 => x"3482b6a4",
          2553 => x"088c0508",
          2554 => x"5380730c",
          2555 => x"82b6a408",
          2556 => x"88050870",
          2557 => x"08515372",
          2558 => x"33537282",
          2559 => x"b6a408f8",
          2560 => x"05347281",
          2561 => x"ff065372",
          2562 => x"a02e0981",
          2563 => x"06913882",
          2564 => x"b6a40888",
          2565 => x"05087008",
          2566 => x"8105710c",
          2567 => x"53ce3982",
          2568 => x"b6a408f8",
          2569 => x"05335372",
          2570 => x"ad2e0981",
          2571 => x"06a43881",
          2572 => x"0b82b6a4",
          2573 => x"08f00534",
          2574 => x"82b6a408",
          2575 => x"88050870",
          2576 => x"08810571",
          2577 => x"0c700851",
          2578 => x"53723382",
          2579 => x"b6a408f8",
          2580 => x"053482b6",
          2581 => x"a408f805",
          2582 => x"335372b0",
          2583 => x"2e098106",
          2584 => x"81dc3882",
          2585 => x"b6a40888",
          2586 => x"05087008",
          2587 => x"8105710c",
          2588 => x"70085153",
          2589 => x"723382b6",
          2590 => x"a408f805",
          2591 => x"3482b6a4",
          2592 => x"08f80533",
          2593 => x"82b6a408",
          2594 => x"e8050c82",
          2595 => x"b6a408e8",
          2596 => x"050880e2",
          2597 => x"2eb63882",
          2598 => x"b6a408e8",
          2599 => x"050880f8",
          2600 => x"2e843880",
          2601 => x"cd39900b",
          2602 => x"82b6a408",
          2603 => x"f4053482",
          2604 => x"b6a40888",
          2605 => x"05087008",
          2606 => x"8105710c",
          2607 => x"70085153",
          2608 => x"723382b6",
          2609 => x"a408f805",
          2610 => x"3481a439",
          2611 => x"820b82b6",
          2612 => x"a408f405",
          2613 => x"3482b6a4",
          2614 => x"08880508",
          2615 => x"70088105",
          2616 => x"710c7008",
          2617 => x"51537233",
          2618 => x"82b6a408",
          2619 => x"f8053480",
          2620 => x"fe3982b6",
          2621 => x"a408f805",
          2622 => x"335372a0",
          2623 => x"268d3881",
          2624 => x"0b82b6a4",
          2625 => x"08ec050c",
          2626 => x"83803982",
          2627 => x"b6a408f8",
          2628 => x"053353af",
          2629 => x"73279038",
          2630 => x"82b6a408",
          2631 => x"f8053353",
          2632 => x"72b92683",
          2633 => x"388d3980",
          2634 => x"0b82b6a4",
          2635 => x"08ec050c",
          2636 => x"82d83988",
          2637 => x"0b82b6a4",
          2638 => x"08f40534",
          2639 => x"b23982b6",
          2640 => x"a408f805",
          2641 => x"3353af73",
          2642 => x"27903882",
          2643 => x"b6a408f8",
          2644 => x"05335372",
          2645 => x"b9268338",
          2646 => x"8d39800b",
          2647 => x"82b6a408",
          2648 => x"ec050c82",
          2649 => x"a5398a0b",
          2650 => x"82b6a408",
          2651 => x"f4053480",
          2652 => x"0b82b6a4",
          2653 => x"08fc050c",
          2654 => x"82b6a408",
          2655 => x"f8053353",
          2656 => x"a0732781",
          2657 => x"cf3882b6",
          2658 => x"a408f805",
          2659 => x"335380e0",
          2660 => x"73279438",
          2661 => x"82b6a408",
          2662 => x"f80533e0",
          2663 => x"11515372",
          2664 => x"82b6a408",
          2665 => x"f8053482",
          2666 => x"b6a408f8",
          2667 => x"0533d011",
          2668 => x"51537282",
          2669 => x"b6a408f8",
          2670 => x"053482b6",
          2671 => x"a408f805",
          2672 => x"33539073",
          2673 => x"27ad3882",
          2674 => x"b6a408f8",
          2675 => x"0533f911",
          2676 => x"51537282",
          2677 => x"b6a408f8",
          2678 => x"053482b6",
          2679 => x"a408f805",
          2680 => x"33537289",
          2681 => x"268d3880",
          2682 => x"0b82b6a4",
          2683 => x"08ec050c",
          2684 => x"81983982",
          2685 => x"b6a408f8",
          2686 => x"053382b6",
          2687 => x"a408f405",
          2688 => x"33545472",
          2689 => x"74268d38",
          2690 => x"800b82b6",
          2691 => x"a408ec05",
          2692 => x"0c80f739",
          2693 => x"82b6a408",
          2694 => x"f4053370",
          2695 => x"82b6a408",
          2696 => x"fc050829",
          2697 => x"82b6a408",
          2698 => x"f8053370",
          2699 => x"1282b6a4",
          2700 => x"08fc050c",
          2701 => x"82b6a408",
          2702 => x"88050870",
          2703 => x"08810571",
          2704 => x"0c700851",
          2705 => x"51525553",
          2706 => x"723382b6",
          2707 => x"a408f805",
          2708 => x"34fea539",
          2709 => x"82b6a408",
          2710 => x"f0053353",
          2711 => x"72802e90",
          2712 => x"3882b6a4",
          2713 => x"08fc0508",
          2714 => x"3082b6a4",
          2715 => x"08fc050c",
          2716 => x"82b6a408",
          2717 => x"8c050882",
          2718 => x"b6a408fc",
          2719 => x"0508710c",
          2720 => x"53810b82",
          2721 => x"b6a408ec",
          2722 => x"050c82b6",
          2723 => x"a408ec05",
          2724 => x"0882b698",
          2725 => x"0c8b3d0d",
          2726 => x"82b6a40c",
          2727 => x"04f93d0d",
          2728 => x"79700870",
          2729 => x"56565874",
          2730 => x"802e80e3",
          2731 => x"38953975",
          2732 => x"0851e6d1",
          2733 => x"3f82b698",
          2734 => x"0815780c",
          2735 => x"85163354",
          2736 => x"80cd3974",
          2737 => x"335473a0",
          2738 => x"2e098106",
          2739 => x"86388115",
          2740 => x"55f13980",
          2741 => x"57769029",
          2742 => x"82b19805",
          2743 => x"70085256",
          2744 => x"e6a33f82",
          2745 => x"b6980853",
          2746 => x"74527508",
          2747 => x"51e9a33f",
          2748 => x"82b69808",
          2749 => x"8b388416",
          2750 => x"33547381",
          2751 => x"2effb038",
          2752 => x"81177081",
          2753 => x"ff065854",
          2754 => x"997727c9",
          2755 => x"38ff5473",
          2756 => x"82b6980c",
          2757 => x"893d0d04",
          2758 => x"ff3d0d73",
          2759 => x"52719326",
          2760 => x"818e3871",
          2761 => x"84298295",
          2762 => x"cc055271",
          2763 => x"0804829b",
          2764 => x"98518180",
          2765 => x"39829ba4",
          2766 => x"5180f939",
          2767 => x"829bb451",
          2768 => x"80f23982",
          2769 => x"9bc45180",
          2770 => x"eb39829b",
          2771 => x"d45180e4",
          2772 => x"39829be4",
          2773 => x"5180dd39",
          2774 => x"829bf851",
          2775 => x"80d63982",
          2776 => x"9c885180",
          2777 => x"cf39829c",
          2778 => x"a05180c8",
          2779 => x"39829cb8",
          2780 => x"5180c139",
          2781 => x"829cd051",
          2782 => x"bb39829c",
          2783 => x"ec51b539",
          2784 => x"829d8051",
          2785 => x"af39829d",
          2786 => x"a851a939",
          2787 => x"829db851",
          2788 => x"a339829d",
          2789 => x"d8519d39",
          2790 => x"829de851",
          2791 => x"9739829e",
          2792 => x"80519139",
          2793 => x"829e9851",
          2794 => x"8b39829e",
          2795 => x"b0518539",
          2796 => x"829ebc51",
          2797 => x"d8ad3f83",
          2798 => x"3d0d04fb",
          2799 => x"3d0d7779",
          2800 => x"56567487",
          2801 => x"e7268a38",
          2802 => x"74527587",
          2803 => x"e8295190",
          2804 => x"3987e852",
          2805 => x"7451efab",
          2806 => x"3f82b698",
          2807 => x"08527551",
          2808 => x"efa13f82",
          2809 => x"b6980854",
          2810 => x"79537552",
          2811 => x"829ecc51",
          2812 => x"ffbbe53f",
          2813 => x"873d0d04",
          2814 => x"ec3d0d66",
          2815 => x"02840580",
          2816 => x"e305335b",
          2817 => x"57806878",
          2818 => x"30707a07",
          2819 => x"73255157",
          2820 => x"59597856",
          2821 => x"7787ff26",
          2822 => x"83388156",
          2823 => x"74760770",
          2824 => x"81ff0651",
          2825 => x"55935674",
          2826 => x"81823881",
          2827 => x"5376528c",
          2828 => x"3d705256",
          2829 => x"80ffe73f",
          2830 => x"82b69808",
          2831 => x"5782b698",
          2832 => x"08b93882",
          2833 => x"b6980887",
          2834 => x"c098880c",
          2835 => x"82b69808",
          2836 => x"59963dd4",
          2837 => x"05548480",
          2838 => x"53775275",
          2839 => x"518184a3",
          2840 => x"3f82b698",
          2841 => x"085782b6",
          2842 => x"98089038",
          2843 => x"7a557480",
          2844 => x"2e893874",
          2845 => x"19751959",
          2846 => x"59d73996",
          2847 => x"3dd80551",
          2848 => x"818c8c3f",
          2849 => x"76307078",
          2850 => x"0780257b",
          2851 => x"30709f2a",
          2852 => x"72065157",
          2853 => x"51567480",
          2854 => x"2e903882",
          2855 => x"9ef05387",
          2856 => x"c0988808",
          2857 => x"527851fe",
          2858 => x"923f7656",
          2859 => x"7582b698",
          2860 => x"0c963d0d",
          2861 => x"04f73d0d",
          2862 => x"7d028405",
          2863 => x"bb053359",
          2864 => x"5aff5980",
          2865 => x"537c527b",
          2866 => x"51fead3f",
          2867 => x"82b69808",
          2868 => x"80cb3877",
          2869 => x"802e8838",
          2870 => x"77812ebf",
          2871 => x"38bf3982",
          2872 => x"cde85782",
          2873 => x"cde85682",
          2874 => x"cde85582",
          2875 => x"cdf00854",
          2876 => x"82cdec08",
          2877 => x"5382cde8",
          2878 => x"0852829e",
          2879 => x"f851ffb9",
          2880 => x"d73f82cd",
          2881 => x"e8566255",
          2882 => x"615482b6",
          2883 => x"98536052",
          2884 => x"7f51792d",
          2885 => x"82b69808",
          2886 => x"59833979",
          2887 => x"047882b6",
          2888 => x"980c8b3d",
          2889 => x"0d04f33d",
          2890 => x"0d7f6163",
          2891 => x"028c0580",
          2892 => x"cf053373",
          2893 => x"73156841",
          2894 => x"5f5c5c5e",
          2895 => x"5e5e7a52",
          2896 => x"829fac51",
          2897 => x"ffb9913f",
          2898 => x"829fb451",
          2899 => x"ffb9893f",
          2900 => x"80557479",
          2901 => x"27818038",
          2902 => x"7b902e89",
          2903 => x"387ba02e",
          2904 => x"a73880c6",
          2905 => x"39741853",
          2906 => x"727a278e",
          2907 => x"38722252",
          2908 => x"829fb851",
          2909 => x"ffb8e13f",
          2910 => x"8939829f",
          2911 => x"c451ffb8",
          2912 => x"d73f8215",
          2913 => x"5580c339",
          2914 => x"74185372",
          2915 => x"7a278e38",
          2916 => x"72085282",
          2917 => x"9fac51ff",
          2918 => x"b8be3f89",
          2919 => x"39829fc0",
          2920 => x"51ffb8b4",
          2921 => x"3f841555",
          2922 => x"a1397418",
          2923 => x"53727a27",
          2924 => x"8e387233",
          2925 => x"52829fcc",
          2926 => x"51ffb89c",
          2927 => x"3f893982",
          2928 => x"9fd451ff",
          2929 => x"b8923f81",
          2930 => x"155582cd",
          2931 => x"ec0852a0",
          2932 => x"51d7df3f",
          2933 => x"fefc3982",
          2934 => x"9fd851ff",
          2935 => x"b7fa3f80",
          2936 => x"55747927",
          2937 => x"80c63874",
          2938 => x"18703355",
          2939 => x"53805672",
          2940 => x"7a278338",
          2941 => x"81568053",
          2942 => x"9f742783",
          2943 => x"38815375",
          2944 => x"73067081",
          2945 => x"ff065153",
          2946 => x"72802e90",
          2947 => x"387380fe",
          2948 => x"268a3882",
          2949 => x"cdec0852",
          2950 => x"73518839",
          2951 => x"82cdec08",
          2952 => x"52a051d7",
          2953 => x"8d3f8115",
          2954 => x"55ffb639",
          2955 => x"829fdc51",
          2956 => x"d3b13f78",
          2957 => x"18791c5c",
          2958 => x"589ccb3f",
          2959 => x"82b69808",
          2960 => x"982b7098",
          2961 => x"2c515776",
          2962 => x"a02e0981",
          2963 => x"06aa389c",
          2964 => x"b53f82b6",
          2965 => x"9808982b",
          2966 => x"70982c70",
          2967 => x"a0327030",
          2968 => x"729b3270",
          2969 => x"30707207",
          2970 => x"73750706",
          2971 => x"51585859",
          2972 => x"57515780",
          2973 => x"7324d838",
          2974 => x"769b2e09",
          2975 => x"81068538",
          2976 => x"80538c39",
          2977 => x"7c1e5372",
          2978 => x"7826fdb2",
          2979 => x"38ff5372",
          2980 => x"82b6980c",
          2981 => x"8f3d0d04",
          2982 => x"fc3d0d02",
          2983 => x"9b053382",
          2984 => x"9fe05382",
          2985 => x"9fe45255",
          2986 => x"ffb6ad3f",
          2987 => x"82b4f022",
          2988 => x"51a5a43f",
          2989 => x"829ff054",
          2990 => x"829ffc53",
          2991 => x"82b4f133",
          2992 => x"5282a084",
          2993 => x"51ffb690",
          2994 => x"3f74802e",
          2995 => x"8438a0d8",
          2996 => x"3f863d0d",
          2997 => x"04fe3d0d",
          2998 => x"87c09680",
          2999 => x"0853a5c0",
          3000 => x"3f815198",
          3001 => x"8e3f82a0",
          3002 => x"a05199a3",
          3003 => x"3f805198",
          3004 => x"823f7281",
          3005 => x"2a708106",
          3006 => x"51527180",
          3007 => x"2e923881",
          3008 => x"5197f03f",
          3009 => x"82a0b851",
          3010 => x"99853f80",
          3011 => x"5197e43f",
          3012 => x"72822a70",
          3013 => x"81065152",
          3014 => x"71802e92",
          3015 => x"38815197",
          3016 => x"d23f82a0",
          3017 => x"c85198e7",
          3018 => x"3f805197",
          3019 => x"c63f7283",
          3020 => x"2a708106",
          3021 => x"51527180",
          3022 => x"2e923881",
          3023 => x"5197b43f",
          3024 => x"82a0d851",
          3025 => x"98c93f80",
          3026 => x"5197a83f",
          3027 => x"72842a70",
          3028 => x"81065152",
          3029 => x"71802e92",
          3030 => x"38815197",
          3031 => x"963f82a0",
          3032 => x"ec5198ab",
          3033 => x"3f805197",
          3034 => x"8a3f7285",
          3035 => x"2a708106",
          3036 => x"51527180",
          3037 => x"2e923881",
          3038 => x"5196f83f",
          3039 => x"82a18051",
          3040 => x"988d3f80",
          3041 => x"5196ec3f",
          3042 => x"72862a70",
          3043 => x"81065152",
          3044 => x"71802e92",
          3045 => x"38815196",
          3046 => x"da3f82a1",
          3047 => x"945197ef",
          3048 => x"3f805196",
          3049 => x"ce3f7287",
          3050 => x"2a708106",
          3051 => x"51527180",
          3052 => x"2e923881",
          3053 => x"5196bc3f",
          3054 => x"82a1a851",
          3055 => x"97d13f80",
          3056 => x"5196b03f",
          3057 => x"72882a70",
          3058 => x"81065152",
          3059 => x"71802e92",
          3060 => x"38815196",
          3061 => x"9e3f82a1",
          3062 => x"bc5197b3",
          3063 => x"3f805196",
          3064 => x"923fa3c4",
          3065 => x"3f843d0d",
          3066 => x"04fb3d0d",
          3067 => x"77028405",
          3068 => x"a3053370",
          3069 => x"55565680",
          3070 => x"527551e2",
          3071 => x"e93f0b0b",
          3072 => x"82b19433",
          3073 => x"5473a938",
          3074 => x"815382a1",
          3075 => x"f85282cd",
          3076 => x"985180f8",
          3077 => x"893f82b6",
          3078 => x"98083070",
          3079 => x"82b69808",
          3080 => x"07802582",
          3081 => x"71315151",
          3082 => x"54730b0b",
          3083 => x"82b19434",
          3084 => x"0b0b82b1",
          3085 => x"94335473",
          3086 => x"812e0981",
          3087 => x"06af3882",
          3088 => x"cd985374",
          3089 => x"52755181",
          3090 => x"b2ba3f82",
          3091 => x"b6980880",
          3092 => x"2e8b3882",
          3093 => x"b6980851",
          3094 => x"cf893f91",
          3095 => x"3982cd98",
          3096 => x"518184ab",
          3097 => x"3f820b0b",
          3098 => x"0b82b194",
          3099 => x"340b0b82",
          3100 => x"b1943354",
          3101 => x"73822e09",
          3102 => x"81068c38",
          3103 => x"82a28853",
          3104 => x"74527551",
          3105 => x"a9bc3f80",
          3106 => x"0b82b698",
          3107 => x"0c873d0d",
          3108 => x"04ce3d0d",
          3109 => x"80707182",
          3110 => x"cd940c5f",
          3111 => x"5d81527c",
          3112 => x"5180c6d5",
          3113 => x"3f82b698",
          3114 => x"0881ff06",
          3115 => x"59787d2e",
          3116 => x"098106a3",
          3117 => x"38963d59",
          3118 => x"835382a2",
          3119 => x"90527851",
          3120 => x"dca33f7c",
          3121 => x"53785282",
          3122 => x"b7c45180",
          3123 => x"f5ef3f82",
          3124 => x"b698087d",
          3125 => x"2e883882",
          3126 => x"a294518d",
          3127 => x"a3398170",
          3128 => x"5f5d82a2",
          3129 => x"cc51ffb1",
          3130 => x"ef3f963d",
          3131 => x"70465a80",
          3132 => x"f8527951",
          3133 => x"fdf33fb4",
          3134 => x"3dff8405",
          3135 => x"51f39e3f",
          3136 => x"82b69808",
          3137 => x"902b7090",
          3138 => x"2c515978",
          3139 => x"80c22e87",
          3140 => x"a3387880",
          3141 => x"c224b238",
          3142 => x"78bd2e81",
          3143 => x"d23878bd",
          3144 => x"24903878",
          3145 => x"802effba",
          3146 => x"3878bc2e",
          3147 => x"80da388a",
          3148 => x"d4397880",
          3149 => x"c02e8399",
          3150 => x"387880c0",
          3151 => x"2485cd38",
          3152 => x"78bf2e82",
          3153 => x"8c388abd",
          3154 => x"397880f9",
          3155 => x"2e89d938",
          3156 => x"7880f924",
          3157 => x"92387880",
          3158 => x"c32e8888",
          3159 => x"387880f8",
          3160 => x"2e89a138",
          3161 => x"8a9f3978",
          3162 => x"81832e8a",
          3163 => x"86387881",
          3164 => x"83248b38",
          3165 => x"7881822e",
          3166 => x"89eb388a",
          3167 => x"88397881",
          3168 => x"852e89fb",
          3169 => x"3889fe39",
          3170 => x"b43dff80",
          3171 => x"1153ff84",
          3172 => x"0551ecb8",
          3173 => x"3f82b698",
          3174 => x"08802efe",
          3175 => x"c538b43d",
          3176 => x"fefc1153",
          3177 => x"ff840551",
          3178 => x"eca23f82",
          3179 => x"b6980880",
          3180 => x"2efeaf38",
          3181 => x"b43dfef8",
          3182 => x"1153ff84",
          3183 => x"0551ec8c",
          3184 => x"3f82b698",
          3185 => x"08863882",
          3186 => x"b6980842",
          3187 => x"82a2d051",
          3188 => x"ffb0853f",
          3189 => x"63635c5a",
          3190 => x"797b2781",
          3191 => x"ec386159",
          3192 => x"787a7084",
          3193 => x"055c0c7a",
          3194 => x"7a26f538",
          3195 => x"81db39b4",
          3196 => x"3dff8011",
          3197 => x"53ff8405",
          3198 => x"51ebd13f",
          3199 => x"82b69808",
          3200 => x"802efdde",
          3201 => x"38b43dfe",
          3202 => x"fc1153ff",
          3203 => x"840551eb",
          3204 => x"bb3f82b6",
          3205 => x"9808802e",
          3206 => x"fdc838b4",
          3207 => x"3dfef811",
          3208 => x"53ff8405",
          3209 => x"51eba53f",
          3210 => x"82b69808",
          3211 => x"802efdb2",
          3212 => x"3882a2e0",
          3213 => x"51ffafa0",
          3214 => x"3f635a79",
          3215 => x"63278189",
          3216 => x"38615979",
          3217 => x"7081055b",
          3218 => x"33793461",
          3219 => x"810542eb",
          3220 => x"39b43dff",
          3221 => x"801153ff",
          3222 => x"840551ea",
          3223 => x"ef3f82b6",
          3224 => x"9808802e",
          3225 => x"fcfc38b4",
          3226 => x"3dfefc11",
          3227 => x"53ff8405",
          3228 => x"51ead93f",
          3229 => x"82b69808",
          3230 => x"802efce6",
          3231 => x"38b43dfe",
          3232 => x"f81153ff",
          3233 => x"840551ea",
          3234 => x"c33f82b6",
          3235 => x"9808802e",
          3236 => x"fcd03882",
          3237 => x"a2ec51ff",
          3238 => x"aebe3f63",
          3239 => x"5a796327",
          3240 => x"a8386170",
          3241 => x"337b335e",
          3242 => x"5a5b787c",
          3243 => x"2e923878",
          3244 => x"557a5479",
          3245 => x"33537952",
          3246 => x"82a2fc51",
          3247 => x"ffae993f",
          3248 => x"811a6281",
          3249 => x"05435ad5",
          3250 => x"398a51cd",
          3251 => x"b83ffc92",
          3252 => x"39b43dff",
          3253 => x"801153ff",
          3254 => x"840551e9",
          3255 => x"ef3f82b6",
          3256 => x"980880df",
          3257 => x"3882b584",
          3258 => x"33597880",
          3259 => x"2e893882",
          3260 => x"b4bc0844",
          3261 => x"80cd3982",
          3262 => x"b5853359",
          3263 => x"78802e88",
          3264 => x"3882b4c4",
          3265 => x"0844bc39",
          3266 => x"82b58633",
          3267 => x"5978802e",
          3268 => x"883882b4",
          3269 => x"cc0844ab",
          3270 => x"3982b587",
          3271 => x"33597880",
          3272 => x"2e883882",
          3273 => x"b4d40844",
          3274 => x"9a3982b5",
          3275 => x"82335978",
          3276 => x"802e8838",
          3277 => x"82b4dc08",
          3278 => x"44893982",
          3279 => x"b4ec08fc",
          3280 => x"800544b4",
          3281 => x"3dfefc11",
          3282 => x"53ff8405",
          3283 => x"51e8fd3f",
          3284 => x"82b69808",
          3285 => x"80de3882",
          3286 => x"b5843359",
          3287 => x"78802e89",
          3288 => x"3882b4c0",
          3289 => x"084380cc",
          3290 => x"3982b585",
          3291 => x"33597880",
          3292 => x"2e883882",
          3293 => x"b4c80843",
          3294 => x"bb3982b5",
          3295 => x"86335978",
          3296 => x"802e8838",
          3297 => x"82b4d008",
          3298 => x"43aa3982",
          3299 => x"b5873359",
          3300 => x"78802e88",
          3301 => x"3882b4d8",
          3302 => x"08439939",
          3303 => x"82b58233",
          3304 => x"5978802e",
          3305 => x"883882b4",
          3306 => x"e0084388",
          3307 => x"3982b4ec",
          3308 => x"08880543",
          3309 => x"b43dfef8",
          3310 => x"1153ff84",
          3311 => x"0551e88c",
          3312 => x"3f82b698",
          3313 => x"08802ea7",
          3314 => x"3880625c",
          3315 => x"5c7a882e",
          3316 => x"8338815c",
          3317 => x"7a903270",
          3318 => x"30707207",
          3319 => x"9f2a707f",
          3320 => x"0651515a",
          3321 => x"5a78802e",
          3322 => x"88387aa0",
          3323 => x"2e833888",
          3324 => x"4282a398",
          3325 => x"51c7ec3f",
          3326 => x"a0556354",
          3327 => x"61536252",
          3328 => x"6351f2a2",
          3329 => x"3f82a3a4",
          3330 => x"5186f539",
          3331 => x"b43dff80",
          3332 => x"1153ff84",
          3333 => x"0551e7b4",
          3334 => x"3f82b698",
          3335 => x"08802ef9",
          3336 => x"c138b43d",
          3337 => x"fefc1153",
          3338 => x"ff840551",
          3339 => x"e79e3f82",
          3340 => x"b6980880",
          3341 => x"2ea43863",
          3342 => x"590280cb",
          3343 => x"05337934",
          3344 => x"63810544",
          3345 => x"b43dfefc",
          3346 => x"1153ff84",
          3347 => x"0551e6fc",
          3348 => x"3f82b698",
          3349 => x"08e138f9",
          3350 => x"89396370",
          3351 => x"33545282",
          3352 => x"a3b051ff",
          3353 => x"aaf23f82",
          3354 => x"cde80853",
          3355 => x"80f85279",
          3356 => x"51ffabb9",
          3357 => x"3f794579",
          3358 => x"335978ae",
          3359 => x"2ef8e338",
          3360 => x"9f79279f",
          3361 => x"38b43dfe",
          3362 => x"fc1153ff",
          3363 => x"840551e6",
          3364 => x"bb3f82b6",
          3365 => x"9808802e",
          3366 => x"91386359",
          3367 => x"0280cb05",
          3368 => x"33793463",
          3369 => x"810544ff",
          3370 => x"b13982a3",
          3371 => x"bc51c6b3",
          3372 => x"3fffa739",
          3373 => x"b43dfef4",
          3374 => x"1153ff84",
          3375 => x"0551e0bb",
          3376 => x"3f82b698",
          3377 => x"08802ef8",
          3378 => x"9938b43d",
          3379 => x"fef01153",
          3380 => x"ff840551",
          3381 => x"e0a53f82",
          3382 => x"b6980880",
          3383 => x"2ea53860",
          3384 => x"5902be05",
          3385 => x"22797082",
          3386 => x"055b2378",
          3387 => x"41b43dfe",
          3388 => x"f01153ff",
          3389 => x"840551e0",
          3390 => x"823f82b6",
          3391 => x"9808e038",
          3392 => x"f7e03960",
          3393 => x"70225452",
          3394 => x"82a3c051",
          3395 => x"ffa9c93f",
          3396 => x"82cde808",
          3397 => x"5380f852",
          3398 => x"7951ffaa",
          3399 => x"903f7945",
          3400 => x"79335978",
          3401 => x"ae2ef7ba",
          3402 => x"38789f26",
          3403 => x"87386082",
          3404 => x"0541d039",
          3405 => x"b43dfef0",
          3406 => x"1153ff84",
          3407 => x"0551dfbb",
          3408 => x"3f82b698",
          3409 => x"08802e92",
          3410 => x"38605902",
          3411 => x"be052279",
          3412 => x"7082055b",
          3413 => x"237841ff",
          3414 => x"aa3982a3",
          3415 => x"bc51c583",
          3416 => x"3fffa039",
          3417 => x"b43dfef4",
          3418 => x"1153ff84",
          3419 => x"0551df8b",
          3420 => x"3f82b698",
          3421 => x"08802ef6",
          3422 => x"e938b43d",
          3423 => x"fef01153",
          3424 => x"ff840551",
          3425 => x"def53f82",
          3426 => x"b6980880",
          3427 => x"2ea03860",
          3428 => x"60710c59",
          3429 => x"60840541",
          3430 => x"b43dfef0",
          3431 => x"1153ff84",
          3432 => x"0551ded7",
          3433 => x"3f82b698",
          3434 => x"08e538f6",
          3435 => x"b5396070",
          3436 => x"08545282",
          3437 => x"a3cc51ff",
          3438 => x"a89e3f82",
          3439 => x"cde80853",
          3440 => x"80f85279",
          3441 => x"51ffa8e5",
          3442 => x"3f794579",
          3443 => x"335978ae",
          3444 => x"2ef68f38",
          3445 => x"9f79279b",
          3446 => x"38b43dfe",
          3447 => x"f01153ff",
          3448 => x"840551de",
          3449 => x"963f82b6",
          3450 => x"9808802e",
          3451 => x"8d386060",
          3452 => x"710c5960",
          3453 => x"840541ff",
          3454 => x"b53982a3",
          3455 => x"bc51c3e3",
          3456 => x"3fffab39",
          3457 => x"b43dff80",
          3458 => x"1153ff84",
          3459 => x"0551e3bc",
          3460 => x"3f82b698",
          3461 => x"08802ef5",
          3462 => x"c9386352",
          3463 => x"82a3dc51",
          3464 => x"ffa7b53f",
          3465 => x"63597804",
          3466 => x"b43dff80",
          3467 => x"1153ff84",
          3468 => x"0551e398",
          3469 => x"3f82b698",
          3470 => x"08802ef5",
          3471 => x"a5386352",
          3472 => x"82a3f851",
          3473 => x"ffa7913f",
          3474 => x"6359782d",
          3475 => x"82b69808",
          3476 => x"802ef58e",
          3477 => x"3882b698",
          3478 => x"085282a4",
          3479 => x"9451ffa6",
          3480 => x"f73ff4fe",
          3481 => x"3982a4b0",
          3482 => x"51c2f83f",
          3483 => x"ffa6ca3f",
          3484 => x"f4f03982",
          3485 => x"a4cc51c2",
          3486 => x"ea3f8059",
          3487 => x"ffa83991",
          3488 => x"a73ff4de",
          3489 => x"39794579",
          3490 => x"33597880",
          3491 => x"2ef4d338",
          3492 => x"7d7d0659",
          3493 => x"78802e81",
          3494 => x"cf38b43d",
          3495 => x"ff840551",
          3496 => x"83ca3f82",
          3497 => x"b698085c",
          3498 => x"815b7a82",
          3499 => x"2eb2387a",
          3500 => x"82248938",
          3501 => x"7a812e8c",
          3502 => x"3880ca39",
          3503 => x"7a832ead",
          3504 => x"3880c239",
          3505 => x"82a4e056",
          3506 => x"7b5582a4",
          3507 => x"e4548053",
          3508 => x"82a4e852",
          3509 => x"b43dffb0",
          3510 => x"0551ffa8",
          3511 => x"e33fb839",
          3512 => x"7b52b43d",
          3513 => x"ffb00551",
          3514 => x"cf893fab",
          3515 => x"397b5582",
          3516 => x"a4e45480",
          3517 => x"5382a4f8",
          3518 => x"52b43dff",
          3519 => x"b00551ff",
          3520 => x"a8be3f93",
          3521 => x"397b5480",
          3522 => x"5382a584",
          3523 => x"52b43dff",
          3524 => x"b00551ff",
          3525 => x"a8aa3f82",
          3526 => x"b4bc5882",
          3527 => x"b6c85780",
          3528 => x"56645580",
          3529 => x"5482d080",
          3530 => x"5382d080",
          3531 => x"52b43dff",
          3532 => x"b00551eb",
          3533 => x"803f82b6",
          3534 => x"980882b6",
          3535 => x"98080970",
          3536 => x"30707207",
          3537 => x"8025515b",
          3538 => x"5b5f805a",
          3539 => x"7a832683",
          3540 => x"38815a78",
          3541 => x"7a065978",
          3542 => x"802e8d38",
          3543 => x"811b7081",
          3544 => x"ff065c59",
          3545 => x"7afec338",
          3546 => x"7d81327d",
          3547 => x"81320759",
          3548 => x"788a387e",
          3549 => x"ff2e0981",
          3550 => x"06f2e738",
          3551 => x"82a58c51",
          3552 => x"c0e13ff2",
          3553 => x"dd39f53d",
          3554 => x"0d800b82",
          3555 => x"b6c83487",
          3556 => x"c0948c70",
          3557 => x"08545587",
          3558 => x"84805272",
          3559 => x"51d7e43f",
          3560 => x"82b69808",
          3561 => x"902b7508",
          3562 => x"55538784",
          3563 => x"80527351",
          3564 => x"d7d13f72",
          3565 => x"82b69808",
          3566 => x"07750c87",
          3567 => x"c0949c70",
          3568 => x"08545587",
          3569 => x"84805272",
          3570 => x"51d7b83f",
          3571 => x"82b69808",
          3572 => x"902b7508",
          3573 => x"55538784",
          3574 => x"80527351",
          3575 => x"d7a53f72",
          3576 => x"82b69808",
          3577 => x"07750c8c",
          3578 => x"80830b87",
          3579 => x"c094840c",
          3580 => x"8c80830b",
          3581 => x"87c09494",
          3582 => x"0c80f68b",
          3583 => x"5a80f8f7",
          3584 => x"5b830284",
          3585 => x"05990534",
          3586 => x"805c82cd",
          3587 => x"e80b873d",
          3588 => x"7088130c",
          3589 => x"70720c82",
          3590 => x"cdec0c54",
          3591 => x"89be3f92",
          3592 => x"ff3f82a5",
          3593 => x"9c51ffbf",
          3594 => x"ba3f82a5",
          3595 => x"a851ffbf",
          3596 => x"b23f80dd",
          3597 => x"d55192e3",
          3598 => x"3f8151ec",
          3599 => x"db3ff0d1",
          3600 => x"3f8004fe",
          3601 => x"3d0d8052",
          3602 => x"83537188",
          3603 => x"2b5287d8",
          3604 => x"3f82b698",
          3605 => x"0881ff06",
          3606 => x"7207ff14",
          3607 => x"54527280",
          3608 => x"25e83871",
          3609 => x"82b6980c",
          3610 => x"843d0d04",
          3611 => x"fc3d0d76",
          3612 => x"70085455",
          3613 => x"80735254",
          3614 => x"72742e81",
          3615 => x"8a387233",
          3616 => x"5170a02e",
          3617 => x"09810686",
          3618 => x"38811353",
          3619 => x"f1397233",
          3620 => x"5170a22e",
          3621 => x"09810686",
          3622 => x"38811353",
          3623 => x"81547252",
          3624 => x"73812e09",
          3625 => x"81069f38",
          3626 => x"84398112",
          3627 => x"52807233",
          3628 => x"525470a2",
          3629 => x"2e833881",
          3630 => x"5470802e",
          3631 => x"9d3873ea",
          3632 => x"38983981",
          3633 => x"12528072",
          3634 => x"33525470",
          3635 => x"a02e8338",
          3636 => x"81547080",
          3637 => x"2e843873",
          3638 => x"ea388072",
          3639 => x"33525470",
          3640 => x"a02e0981",
          3641 => x"06833881",
          3642 => x"5470a232",
          3643 => x"70307080",
          3644 => x"25760751",
          3645 => x"51517080",
          3646 => x"2e883880",
          3647 => x"72708105",
          3648 => x"54347175",
          3649 => x"0c725170",
          3650 => x"82b6980c",
          3651 => x"863d0d04",
          3652 => x"fc3d0d76",
          3653 => x"53720880",
          3654 => x"2e913886",
          3655 => x"3dfc0552",
          3656 => x"7251d7d7",
          3657 => x"3f82b698",
          3658 => x"08853880",
          3659 => x"53833974",
          3660 => x"537282b6",
          3661 => x"980c863d",
          3662 => x"0d04fc3d",
          3663 => x"0d768211",
          3664 => x"33ff0552",
          3665 => x"53815270",
          3666 => x"8b268198",
          3667 => x"38831333",
          3668 => x"ff055182",
          3669 => x"52709e26",
          3670 => x"818a3884",
          3671 => x"13335183",
          3672 => x"52709726",
          3673 => x"80fe3885",
          3674 => x"13335184",
          3675 => x"5270bb26",
          3676 => x"80f23886",
          3677 => x"13335185",
          3678 => x"5270bb26",
          3679 => x"80e63888",
          3680 => x"13225586",
          3681 => x"527487e7",
          3682 => x"2680d938",
          3683 => x"8a132254",
          3684 => x"87527387",
          3685 => x"e72680cc",
          3686 => x"38810b87",
          3687 => x"c0989c0c",
          3688 => x"722287c0",
          3689 => x"98bc0c82",
          3690 => x"133387c0",
          3691 => x"98b80c83",
          3692 => x"133387c0",
          3693 => x"98b40c84",
          3694 => x"133387c0",
          3695 => x"98b00c85",
          3696 => x"133387c0",
          3697 => x"98ac0c86",
          3698 => x"133387c0",
          3699 => x"98a80c74",
          3700 => x"87c098a4",
          3701 => x"0c7387c0",
          3702 => x"98a00c80",
          3703 => x"0b87c098",
          3704 => x"9c0c8052",
          3705 => x"7182b698",
          3706 => x"0c863d0d",
          3707 => x"04f33d0d",
          3708 => x"7f5b87c0",
          3709 => x"989c5d81",
          3710 => x"7d0c87c0",
          3711 => x"98bc085e",
          3712 => x"7d7b2387",
          3713 => x"c098b808",
          3714 => x"5a79821c",
          3715 => x"3487c098",
          3716 => x"b4085a79",
          3717 => x"831c3487",
          3718 => x"c098b008",
          3719 => x"5a79841c",
          3720 => x"3487c098",
          3721 => x"ac085a79",
          3722 => x"851c3487",
          3723 => x"c098a808",
          3724 => x"5a79861c",
          3725 => x"3487c098",
          3726 => x"a4085c7b",
          3727 => x"881c2387",
          3728 => x"c098a008",
          3729 => x"5a798a1c",
          3730 => x"23807d0c",
          3731 => x"7983ffff",
          3732 => x"06597b83",
          3733 => x"ffff0658",
          3734 => x"861b3357",
          3735 => x"851b3356",
          3736 => x"841b3355",
          3737 => x"831b3354",
          3738 => x"821b3353",
          3739 => x"7d83ffff",
          3740 => x"065282a5",
          3741 => x"c051ff9e",
          3742 => x"df3f8f3d",
          3743 => x"0d04fb3d",
          3744 => x"0d029f05",
          3745 => x"3382b4b8",
          3746 => x"337081ff",
          3747 => x"06585555",
          3748 => x"87c09484",
          3749 => x"5175802e",
          3750 => x"863887c0",
          3751 => x"94945170",
          3752 => x"0870962a",
          3753 => x"70810653",
          3754 => x"54527080",
          3755 => x"2e8c3871",
          3756 => x"912a7081",
          3757 => x"06515170",
          3758 => x"d7387281",
          3759 => x"32708106",
          3760 => x"51517080",
          3761 => x"2e8d3871",
          3762 => x"932a7081",
          3763 => x"06515170",
          3764 => x"ffbe3873",
          3765 => x"81ff0651",
          3766 => x"87c09480",
          3767 => x"5270802e",
          3768 => x"863887c0",
          3769 => x"94905274",
          3770 => x"720c7482",
          3771 => x"b6980c87",
          3772 => x"3d0d04ff",
          3773 => x"3d0d028f",
          3774 => x"05337030",
          3775 => x"709f2a51",
          3776 => x"52527082",
          3777 => x"b4b83483",
          3778 => x"3d0d04f9",
          3779 => x"3d0d02a7",
          3780 => x"05335877",
          3781 => x"8a2e0981",
          3782 => x"0687387a",
          3783 => x"528d51eb",
          3784 => x"3f82b4b8",
          3785 => x"337081ff",
          3786 => x"06585687",
          3787 => x"c0948453",
          3788 => x"76802e86",
          3789 => x"3887c094",
          3790 => x"94537208",
          3791 => x"70962a70",
          3792 => x"81065556",
          3793 => x"5472802e",
          3794 => x"8c387391",
          3795 => x"2a708106",
          3796 => x"515372d7",
          3797 => x"38748132",
          3798 => x"70810651",
          3799 => x"5372802e",
          3800 => x"8d387393",
          3801 => x"2a708106",
          3802 => x"515372ff",
          3803 => x"be387581",
          3804 => x"ff065387",
          3805 => x"c0948054",
          3806 => x"72802e86",
          3807 => x"3887c094",
          3808 => x"90547774",
          3809 => x"0c800b82",
          3810 => x"b6980c89",
          3811 => x"3d0d04f9",
          3812 => x"3d0d7954",
          3813 => x"80743370",
          3814 => x"81ff0653",
          3815 => x"53577077",
          3816 => x"2e80fc38",
          3817 => x"7181ff06",
          3818 => x"811582b4",
          3819 => x"b8337081",
          3820 => x"ff065957",
          3821 => x"555887c0",
          3822 => x"94845175",
          3823 => x"802e8638",
          3824 => x"87c09494",
          3825 => x"51700870",
          3826 => x"962a7081",
          3827 => x"06535452",
          3828 => x"70802e8c",
          3829 => x"3871912a",
          3830 => x"70810651",
          3831 => x"5170d738",
          3832 => x"72813270",
          3833 => x"81065151",
          3834 => x"70802e8d",
          3835 => x"3871932a",
          3836 => x"70810651",
          3837 => x"5170ffbe",
          3838 => x"387481ff",
          3839 => x"065187c0",
          3840 => x"94805270",
          3841 => x"802e8638",
          3842 => x"87c09490",
          3843 => x"5277720c",
          3844 => x"81177433",
          3845 => x"7081ff06",
          3846 => x"53535770",
          3847 => x"ff863876",
          3848 => x"82b6980c",
          3849 => x"893d0d04",
          3850 => x"fe3d0d82",
          3851 => x"b4b83370",
          3852 => x"81ff0654",
          3853 => x"5287c094",
          3854 => x"84517280",
          3855 => x"2e863887",
          3856 => x"c0949451",
          3857 => x"70087082",
          3858 => x"2a708106",
          3859 => x"51515170",
          3860 => x"802ee238",
          3861 => x"7181ff06",
          3862 => x"5187c094",
          3863 => x"80527080",
          3864 => x"2e863887",
          3865 => x"c0949052",
          3866 => x"71087081",
          3867 => x"ff0682b6",
          3868 => x"980c5184",
          3869 => x"3d0d04ff",
          3870 => x"af3f82b6",
          3871 => x"980881ff",
          3872 => x"0682b698",
          3873 => x"0c04fe3d",
          3874 => x"0d82b4b8",
          3875 => x"337081ff",
          3876 => x"06525387",
          3877 => x"c0948452",
          3878 => x"70802e86",
          3879 => x"3887c094",
          3880 => x"94527108",
          3881 => x"70822a70",
          3882 => x"81065151",
          3883 => x"51ff5270",
          3884 => x"802ea038",
          3885 => x"7281ff06",
          3886 => x"5187c094",
          3887 => x"80527080",
          3888 => x"2e863887",
          3889 => x"c0949052",
          3890 => x"71087098",
          3891 => x"2b70982c",
          3892 => x"51535171",
          3893 => x"82b6980c",
          3894 => x"843d0d04",
          3895 => x"ff3d0d87",
          3896 => x"c09e8008",
          3897 => x"709c2a8a",
          3898 => x"06515170",
          3899 => x"802e84b4",
          3900 => x"3887c09e",
          3901 => x"a40882b4",
          3902 => x"bc0c87c0",
          3903 => x"9ea80882",
          3904 => x"b4c00c87",
          3905 => x"c09e9408",
          3906 => x"82b4c40c",
          3907 => x"87c09e98",
          3908 => x"0882b4c8",
          3909 => x"0c87c09e",
          3910 => x"9c0882b4",
          3911 => x"cc0c87c0",
          3912 => x"9ea00882",
          3913 => x"b4d00c87",
          3914 => x"c09eac08",
          3915 => x"82b4d40c",
          3916 => x"87c09eb0",
          3917 => x"0882b4d8",
          3918 => x"0c87c09e",
          3919 => x"b40882b4",
          3920 => x"dc0c87c0",
          3921 => x"9eb80882",
          3922 => x"b4e00c87",
          3923 => x"c09ebc08",
          3924 => x"82b4e40c",
          3925 => x"87c09ec0",
          3926 => x"0882b4e8",
          3927 => x"0c87c09e",
          3928 => x"c40882b4",
          3929 => x"ec0c87c0",
          3930 => x"9e800851",
          3931 => x"7082b4f0",
          3932 => x"2387c09e",
          3933 => x"840882b4",
          3934 => x"f40c87c0",
          3935 => x"9e880882",
          3936 => x"b4f80c87",
          3937 => x"c09e8c08",
          3938 => x"82b4fc0c",
          3939 => x"810b82b5",
          3940 => x"8034800b",
          3941 => x"87c09e90",
          3942 => x"08708480",
          3943 => x"0a065152",
          3944 => x"5270802e",
          3945 => x"83388152",
          3946 => x"7182b581",
          3947 => x"34800b87",
          3948 => x"c09e9008",
          3949 => x"7088800a",
          3950 => x"06515252",
          3951 => x"70802e83",
          3952 => x"38815271",
          3953 => x"82b58234",
          3954 => x"800b87c0",
          3955 => x"9e900870",
          3956 => x"90800a06",
          3957 => x"51525270",
          3958 => x"802e8338",
          3959 => x"81527182",
          3960 => x"b5833480",
          3961 => x"0b87c09e",
          3962 => x"90087088",
          3963 => x"80800651",
          3964 => x"52527080",
          3965 => x"2e833881",
          3966 => x"527182b5",
          3967 => x"8434800b",
          3968 => x"87c09e90",
          3969 => x"0870a080",
          3970 => x"80065152",
          3971 => x"5270802e",
          3972 => x"83388152",
          3973 => x"7182b585",
          3974 => x"34800b87",
          3975 => x"c09e9008",
          3976 => x"70908080",
          3977 => x"06515252",
          3978 => x"70802e83",
          3979 => x"38815271",
          3980 => x"82b58634",
          3981 => x"800b87c0",
          3982 => x"9e900870",
          3983 => x"84808006",
          3984 => x"51525270",
          3985 => x"802e8338",
          3986 => x"81527182",
          3987 => x"b5873480",
          3988 => x"0b87c09e",
          3989 => x"90087082",
          3990 => x"80800651",
          3991 => x"52527080",
          3992 => x"2e833881",
          3993 => x"527182b5",
          3994 => x"8834800b",
          3995 => x"87c09e90",
          3996 => x"08708180",
          3997 => x"80065152",
          3998 => x"5270802e",
          3999 => x"83388152",
          4000 => x"7182b589",
          4001 => x"34800b87",
          4002 => x"c09e9008",
          4003 => x"7080c080",
          4004 => x"06515252",
          4005 => x"70802e83",
          4006 => x"38815271",
          4007 => x"82b58a34",
          4008 => x"800b87c0",
          4009 => x"9e900870",
          4010 => x"a0800651",
          4011 => x"52527080",
          4012 => x"2e833881",
          4013 => x"527182b5",
          4014 => x"8b3487c0",
          4015 => x"9e900870",
          4016 => x"98800670",
          4017 => x"8a2a5151",
          4018 => x"517082b5",
          4019 => x"8c34800b",
          4020 => x"87c09e90",
          4021 => x"08708480",
          4022 => x"06515252",
          4023 => x"70802e83",
          4024 => x"38815271",
          4025 => x"82b58d34",
          4026 => x"87c09e90",
          4027 => x"087083f0",
          4028 => x"0670842a",
          4029 => x"51515170",
          4030 => x"82b58e34",
          4031 => x"800b87c0",
          4032 => x"9e900870",
          4033 => x"88065152",
          4034 => x"5270802e",
          4035 => x"83388152",
          4036 => x"7182b58f",
          4037 => x"3487c09e",
          4038 => x"90087087",
          4039 => x"06515170",
          4040 => x"82b59034",
          4041 => x"833d0d04",
          4042 => x"fb3d0d82",
          4043 => x"a5d851ff",
          4044 => x"95a63f82",
          4045 => x"b5803354",
          4046 => x"73802e89",
          4047 => x"3882a5ec",
          4048 => x"51ff9594",
          4049 => x"3f82a680",
          4050 => x"51ffb197",
          4051 => x"3f82b582",
          4052 => x"33547380",
          4053 => x"2e943882",
          4054 => x"b4dc0882",
          4055 => x"b4e00811",
          4056 => x"545282a6",
          4057 => x"9851ff94",
          4058 => x"ef3f82b5",
          4059 => x"87335473",
          4060 => x"802e9438",
          4061 => x"82b4d408",
          4062 => x"82b4d808",
          4063 => x"11545282",
          4064 => x"a6b451ff",
          4065 => x"94d23f82",
          4066 => x"b5843354",
          4067 => x"73802e94",
          4068 => x"3882b4bc",
          4069 => x"0882b4c0",
          4070 => x"08115452",
          4071 => x"82a6d051",
          4072 => x"ff94b53f",
          4073 => x"82b58533",
          4074 => x"5473802e",
          4075 => x"943882b4",
          4076 => x"c40882b4",
          4077 => x"c8081154",
          4078 => x"5282a6ec",
          4079 => x"51ff9498",
          4080 => x"3f82b586",
          4081 => x"33547380",
          4082 => x"2e943882",
          4083 => x"b4cc0882",
          4084 => x"b4d00811",
          4085 => x"545282a7",
          4086 => x"8851ff93",
          4087 => x"fb3f82b5",
          4088 => x"8b335473",
          4089 => x"802e8e38",
          4090 => x"82b58c33",
          4091 => x"5282a7a4",
          4092 => x"51ff93e4",
          4093 => x"3f82b58f",
          4094 => x"33547380",
          4095 => x"2e8e3882",
          4096 => x"b5903352",
          4097 => x"82a7c451",
          4098 => x"ff93cd3f",
          4099 => x"82b58d33",
          4100 => x"5473802e",
          4101 => x"8e3882b5",
          4102 => x"8e335282",
          4103 => x"a7e451ff",
          4104 => x"93b63f82",
          4105 => x"b5813354",
          4106 => x"73802e89",
          4107 => x"3882a884",
          4108 => x"51ffafaf",
          4109 => x"3f82b583",
          4110 => x"33547380",
          4111 => x"2e893882",
          4112 => x"a89851ff",
          4113 => x"af9d3f82",
          4114 => x"b5883354",
          4115 => x"73802e89",
          4116 => x"3882a8a4",
          4117 => x"51ffaf8b",
          4118 => x"3f82b589",
          4119 => x"33547380",
          4120 => x"2e893882",
          4121 => x"a8b051ff",
          4122 => x"aef93f82",
          4123 => x"b58a3354",
          4124 => x"73802e89",
          4125 => x"3882a8b8",
          4126 => x"51ffaee7",
          4127 => x"3f82a8c0",
          4128 => x"51ffaedf",
          4129 => x"3f82b4e4",
          4130 => x"085282a8",
          4131 => x"cc51ff92",
          4132 => x"c73f82b4",
          4133 => x"e8085282",
          4134 => x"a8f451ff",
          4135 => x"92ba3f82",
          4136 => x"b4ec0852",
          4137 => x"82a99c51",
          4138 => x"ff92ad3f",
          4139 => x"82a9c451",
          4140 => x"ffaeb03f",
          4141 => x"82b4f022",
          4142 => x"5282a9cc",
          4143 => x"51ff9298",
          4144 => x"3f82b4f4",
          4145 => x"0856bd84",
          4146 => x"c0527551",
          4147 => x"c5b53f82",
          4148 => x"b69808bd",
          4149 => x"84c02976",
          4150 => x"71315454",
          4151 => x"82b69808",
          4152 => x"5282a9f4",
          4153 => x"51ff91f0",
          4154 => x"3f82b587",
          4155 => x"33547380",
          4156 => x"2ea93882",
          4157 => x"b4f80856",
          4158 => x"bd84c052",
          4159 => x"7551c583",
          4160 => x"3f82b698",
          4161 => x"08bd84c0",
          4162 => x"29767131",
          4163 => x"545482b6",
          4164 => x"98085282",
          4165 => x"aaa051ff",
          4166 => x"91be3f82",
          4167 => x"b5823354",
          4168 => x"73802ea9",
          4169 => x"3882b4fc",
          4170 => x"0856bd84",
          4171 => x"c0527551",
          4172 => x"c4d13f82",
          4173 => x"b69808bd",
          4174 => x"84c02976",
          4175 => x"71315454",
          4176 => x"82b69808",
          4177 => x"5282aacc",
          4178 => x"51ff918c",
          4179 => x"3f8a51ff",
          4180 => x"b0b33f87",
          4181 => x"3d0d04fe",
          4182 => x"3d0d0292",
          4183 => x"0533ff05",
          4184 => x"52718426",
          4185 => x"aa387184",
          4186 => x"2982969c",
          4187 => x"05527108",
          4188 => x"0482aaf8",
          4189 => x"519d3982",
          4190 => x"ab805197",
          4191 => x"3982ab88",
          4192 => x"51913982",
          4193 => x"ab90518b",
          4194 => x"3982ab94",
          4195 => x"51853982",
          4196 => x"ab9c51ff",
          4197 => x"90c23f84",
          4198 => x"3d0d0471",
          4199 => x"88800c04",
          4200 => x"800b87c0",
          4201 => x"96840c04",
          4202 => x"82b59408",
          4203 => x"87c09684",
          4204 => x"0c04fd3d",
          4205 => x"0d76982b",
          4206 => x"70982c79",
          4207 => x"982b7098",
          4208 => x"2c721013",
          4209 => x"70822b51",
          4210 => x"53515451",
          4211 => x"51800b82",
          4212 => x"aba81233",
          4213 => x"55537174",
          4214 => x"259c3882",
          4215 => x"aba41108",
          4216 => x"12028405",
          4217 => x"97053371",
          4218 => x"33525252",
          4219 => x"70722e09",
          4220 => x"81068338",
          4221 => x"81537282",
          4222 => x"b6980c85",
          4223 => x"3d0d04fb",
          4224 => x"3d0d7902",
          4225 => x"8405a305",
          4226 => x"33713355",
          4227 => x"56547280",
          4228 => x"2eb13882",
          4229 => x"cdec0852",
          4230 => x"8851ffaf",
          4231 => x"953f82cd",
          4232 => x"ec0852a0",
          4233 => x"51ffaf8a",
          4234 => x"3f82cdec",
          4235 => x"08528851",
          4236 => x"ffaeff3f",
          4237 => x"7333ff05",
          4238 => x"53727434",
          4239 => x"7281ff06",
          4240 => x"53cc3977",
          4241 => x"51ff8f90",
          4242 => x"3f747434",
          4243 => x"873d0d04",
          4244 => x"f63d0d7c",
          4245 => x"028405b7",
          4246 => x"05330288",
          4247 => x"05bb0533",
          4248 => x"82b5f033",
          4249 => x"70842982",
          4250 => x"b5980570",
          4251 => x"08515959",
          4252 => x"5a585974",
          4253 => x"802e8638",
          4254 => x"74519afa",
          4255 => x"3f82b5f0",
          4256 => x"33708429",
          4257 => x"82b59805",
          4258 => x"81197054",
          4259 => x"58565a9d",
          4260 => x"fb3f82b6",
          4261 => x"9808750c",
          4262 => x"82b5f033",
          4263 => x"70842982",
          4264 => x"b5980570",
          4265 => x"0851565a",
          4266 => x"74802ea7",
          4267 => x"38755378",
          4268 => x"527451ff",
          4269 => x"b8af3f82",
          4270 => x"b5f03381",
          4271 => x"05557482",
          4272 => x"b5f03474",
          4273 => x"81ff0655",
          4274 => x"93752787",
          4275 => x"38800b82",
          4276 => x"b5f03477",
          4277 => x"802eb638",
          4278 => x"82b5ec08",
          4279 => x"5675802e",
          4280 => x"ac3882b5",
          4281 => x"e8335574",
          4282 => x"a4388c3d",
          4283 => x"fc055476",
          4284 => x"53785275",
          4285 => x"5180da88",
          4286 => x"3f82b5ec",
          4287 => x"08528a51",
          4288 => x"818f953f",
          4289 => x"82b5ec08",
          4290 => x"5180dde5",
          4291 => x"3f8c3d0d",
          4292 => x"04fd3d0d",
          4293 => x"82b59853",
          4294 => x"93547208",
          4295 => x"5271802e",
          4296 => x"89387151",
          4297 => x"99d03f80",
          4298 => x"730cff14",
          4299 => x"84145454",
          4300 => x"738025e6",
          4301 => x"38800b82",
          4302 => x"b5f03482",
          4303 => x"b5ec0852",
          4304 => x"71802e95",
          4305 => x"38715180",
          4306 => x"dec53f82",
          4307 => x"b5ec0851",
          4308 => x"99a43f80",
          4309 => x"0b82b5ec",
          4310 => x"0c853d0d",
          4311 => x"04dc3d0d",
          4312 => x"81578052",
          4313 => x"82b5ec08",
          4314 => x"5180e3b2",
          4315 => x"3f82b698",
          4316 => x"0880d338",
          4317 => x"82b5ec08",
          4318 => x"5380f852",
          4319 => x"883d7052",
          4320 => x"56818c80",
          4321 => x"3f82b698",
          4322 => x"08802eba",
          4323 => x"387551ff",
          4324 => x"b4f33f82",
          4325 => x"b6980855",
          4326 => x"800b82b6",
          4327 => x"9808259d",
          4328 => x"3882b698",
          4329 => x"08ff0570",
          4330 => x"17555580",
          4331 => x"74347553",
          4332 => x"76528117",
          4333 => x"82ae9852",
          4334 => x"57ff8c9c",
          4335 => x"3f74ff2e",
          4336 => x"098106ff",
          4337 => x"af38a63d",
          4338 => x"0d04d93d",
          4339 => x"0daa3d08",
          4340 => x"ad3d085a",
          4341 => x"5a817058",
          4342 => x"58805282",
          4343 => x"b5ec0851",
          4344 => x"80e2bb3f",
          4345 => x"82b69808",
          4346 => x"819538ff",
          4347 => x"0b82b5ec",
          4348 => x"08545580",
          4349 => x"f8528b3d",
          4350 => x"70525681",
          4351 => x"8b863f82",
          4352 => x"b6980880",
          4353 => x"2ea53875",
          4354 => x"51ffb3f9",
          4355 => x"3f82b698",
          4356 => x"08811858",
          4357 => x"55800b82",
          4358 => x"b6980825",
          4359 => x"8e3882b6",
          4360 => x"9808ff05",
          4361 => x"70175555",
          4362 => x"80743474",
          4363 => x"09703070",
          4364 => x"72079f2a",
          4365 => x"51555578",
          4366 => x"772e8538",
          4367 => x"73ffac38",
          4368 => x"82b5ec08",
          4369 => x"8c110853",
          4370 => x"5180e1d2",
          4371 => x"3f82b698",
          4372 => x"08802e89",
          4373 => x"3882aea4",
          4374 => x"51ff8afc",
          4375 => x"3f78772e",
          4376 => x"0981069b",
          4377 => x"38755279",
          4378 => x"51ffb487",
          4379 => x"3f7951ff",
          4380 => x"b3933fab",
          4381 => x"3d085482",
          4382 => x"b6980874",
          4383 => x"34805877",
          4384 => x"82b6980c",
          4385 => x"a93d0d04",
          4386 => x"f63d0d7c",
          4387 => x"7e715c71",
          4388 => x"72335759",
          4389 => x"5a5873a0",
          4390 => x"2e098106",
          4391 => x"a2387833",
          4392 => x"78055677",
          4393 => x"76279838",
          4394 => x"8117705b",
          4395 => x"70713356",
          4396 => x"585573a0",
          4397 => x"2e098106",
          4398 => x"86387575",
          4399 => x"26ea3880",
          4400 => x"54738829",
          4401 => x"82b5f405",
          4402 => x"70085255",
          4403 => x"ffb2b63f",
          4404 => x"82b69808",
          4405 => x"53795274",
          4406 => x"0851ffb5",
          4407 => x"b53f82b6",
          4408 => x"980880c5",
          4409 => x"38841533",
          4410 => x"5574812e",
          4411 => x"88387482",
          4412 => x"2e8838b5",
          4413 => x"39fce63f",
          4414 => x"ac39811a",
          4415 => x"5a8c3dfc",
          4416 => x"1153f805",
          4417 => x"51c5c53f",
          4418 => x"82b69808",
          4419 => x"802e9a38",
          4420 => x"ff1b5378",
          4421 => x"527751fd",
          4422 => x"b13f82b6",
          4423 => x"980881ff",
          4424 => x"06557485",
          4425 => x"38745491",
          4426 => x"39811470",
          4427 => x"81ff0651",
          4428 => x"54827427",
          4429 => x"ff8b3880",
          4430 => x"547382b6",
          4431 => x"980c8c3d",
          4432 => x"0d04d33d",
          4433 => x"0db03d08",
          4434 => x"b23d08b4",
          4435 => x"3d08595f",
          4436 => x"5a800baf",
          4437 => x"3d3482b5",
          4438 => x"f03382b5",
          4439 => x"ec08555b",
          4440 => x"7381cb38",
          4441 => x"7382b5e8",
          4442 => x"33555573",
          4443 => x"83388155",
          4444 => x"76802e81",
          4445 => x"bc388170",
          4446 => x"76065556",
          4447 => x"73802e81",
          4448 => x"ad38a851",
          4449 => x"98863f82",
          4450 => x"b6980882",
          4451 => x"b5ec0c82",
          4452 => x"b6980880",
          4453 => x"2e819238",
          4454 => x"93537652",
          4455 => x"82b69808",
          4456 => x"5180ccfa",
          4457 => x"3f82b698",
          4458 => x"08802e8c",
          4459 => x"3882aed0",
          4460 => x"51ffa4af",
          4461 => x"3f80f739",
          4462 => x"82b69808",
          4463 => x"5b82b5ec",
          4464 => x"085380f8",
          4465 => x"52903d70",
          4466 => x"52548187",
          4467 => x"b73f82b6",
          4468 => x"98085682",
          4469 => x"b6980874",
          4470 => x"2e098106",
          4471 => x"80d03882",
          4472 => x"b6980851",
          4473 => x"ffb09e3f",
          4474 => x"82b69808",
          4475 => x"55800b82",
          4476 => x"b6980825",
          4477 => x"a93882b6",
          4478 => x"9808ff05",
          4479 => x"70175555",
          4480 => x"80743480",
          4481 => x"537481ff",
          4482 => x"06527551",
          4483 => x"f8c23f81",
          4484 => x"1b7081ff",
          4485 => x"065c5493",
          4486 => x"7b278338",
          4487 => x"805b74ff",
          4488 => x"2e098106",
          4489 => x"ff973886",
          4490 => x"397582b5",
          4491 => x"e834768c",
          4492 => x"3882b5ec",
          4493 => x"08802e84",
          4494 => x"38f9d63f",
          4495 => x"8f3d5dec",
          4496 => x"c53f82b6",
          4497 => x"9808982b",
          4498 => x"70982c51",
          4499 => x"5978ff2e",
          4500 => x"ee387881",
          4501 => x"ff0682cd",
          4502 => x"c4337098",
          4503 => x"2b70982c",
          4504 => x"82cdc033",
          4505 => x"70982b70",
          4506 => x"972c7198",
          4507 => x"2c057084",
          4508 => x"2982aba4",
          4509 => x"05700815",
          4510 => x"70335151",
          4511 => x"51515959",
          4512 => x"51595d58",
          4513 => x"81567378",
          4514 => x"2e80e938",
          4515 => x"777427b4",
          4516 => x"38748180",
          4517 => x"0a2981ff",
          4518 => x"0a057098",
          4519 => x"2c515580",
          4520 => x"752480ce",
          4521 => x"38765374",
          4522 => x"527751f6",
          4523 => x"853f82b6",
          4524 => x"980881ff",
          4525 => x"06547380",
          4526 => x"2ed73874",
          4527 => x"82cdc034",
          4528 => x"8156b139",
          4529 => x"7481800a",
          4530 => x"2981800a",
          4531 => x"0570982c",
          4532 => x"7081ff06",
          4533 => x"56515573",
          4534 => x"95269738",
          4535 => x"76537452",
          4536 => x"7751f5ce",
          4537 => x"3f82b698",
          4538 => x"0881ff06",
          4539 => x"5473cc38",
          4540 => x"d3398056",
          4541 => x"75802e80",
          4542 => x"ca38811c",
          4543 => x"557482cd",
          4544 => x"c4347498",
          4545 => x"2b70982c",
          4546 => x"82cdc033",
          4547 => x"70982b70",
          4548 => x"982c7010",
          4549 => x"1170822b",
          4550 => x"82aba811",
          4551 => x"335e5151",
          4552 => x"51575851",
          4553 => x"5574772e",
          4554 => x"098106fe",
          4555 => x"923882ab",
          4556 => x"ac14087d",
          4557 => x"0c800b82",
          4558 => x"cdc43480",
          4559 => x"0b82cdc0",
          4560 => x"34923975",
          4561 => x"82cdc434",
          4562 => x"7582cdc0",
          4563 => x"3478af3d",
          4564 => x"34757d0c",
          4565 => x"7e547395",
          4566 => x"26fde138",
          4567 => x"73842982",
          4568 => x"96b00554",
          4569 => x"73080482",
          4570 => x"cdcc3354",
          4571 => x"737e2efd",
          4572 => x"cb3882cd",
          4573 => x"c8335573",
          4574 => x"7527ab38",
          4575 => x"74982b70",
          4576 => x"982c5155",
          4577 => x"7375249e",
          4578 => x"38741a54",
          4579 => x"73338115",
          4580 => x"34748180",
          4581 => x"0a2981ff",
          4582 => x"0a057098",
          4583 => x"2c82cdcc",
          4584 => x"33565155",
          4585 => x"df3982cd",
          4586 => x"cc338111",
          4587 => x"56547482",
          4588 => x"cdcc3473",
          4589 => x"1a54ae3d",
          4590 => x"33743482",
          4591 => x"cdc83354",
          4592 => x"737e2589",
          4593 => x"38811454",
          4594 => x"7382cdc8",
          4595 => x"3482cdcc",
          4596 => x"33708180",
          4597 => x"0a2981ff",
          4598 => x"0a057098",
          4599 => x"2c82cdc8",
          4600 => x"335a5156",
          4601 => x"56747725",
          4602 => x"a83882cd",
          4603 => x"ec085274",
          4604 => x"1a703352",
          4605 => x"54ffa3ba",
          4606 => x"3f748180",
          4607 => x"0a298180",
          4608 => x"0a057098",
          4609 => x"2c82cdc8",
          4610 => x"33565155",
          4611 => x"737524da",
          4612 => x"3882cdcc",
          4613 => x"3370982b",
          4614 => x"70982c82",
          4615 => x"cdc8335a",
          4616 => x"51565674",
          4617 => x"7725fc94",
          4618 => x"3882cdec",
          4619 => x"08528851",
          4620 => x"ffa2ff3f",
          4621 => x"7481800a",
          4622 => x"2981800a",
          4623 => x"0570982c",
          4624 => x"82cdc833",
          4625 => x"56515573",
          4626 => x"7524de38",
          4627 => x"fbee3983",
          4628 => x"7a34800b",
          4629 => x"811b3482",
          4630 => x"cdcc5380",
          4631 => x"52829eec",
          4632 => x"51f39c3f",
          4633 => x"81fd3982",
          4634 => x"cdcc3370",
          4635 => x"81ff0655",
          4636 => x"5573802e",
          4637 => x"fbc63882",
          4638 => x"cdc833ff",
          4639 => x"05547382",
          4640 => x"cdc834ff",
          4641 => x"15547382",
          4642 => x"cdcc3482",
          4643 => x"cdec0852",
          4644 => x"8851ffa2",
          4645 => x"9d3f82cd",
          4646 => x"cc337098",
          4647 => x"2b70982c",
          4648 => x"82cdc833",
          4649 => x"57515657",
          4650 => x"747425ad",
          4651 => x"38741a54",
          4652 => x"81143374",
          4653 => x"3482cdec",
          4654 => x"08527333",
          4655 => x"51ffa1f2",
          4656 => x"3f748180",
          4657 => x"0a298180",
          4658 => x"0a057098",
          4659 => x"2c82cdc8",
          4660 => x"33585155",
          4661 => x"757524d5",
          4662 => x"3882cdec",
          4663 => x"0852a051",
          4664 => x"ffa1cf3f",
          4665 => x"82cdcc33",
          4666 => x"70982b70",
          4667 => x"982c82cd",
          4668 => x"c8335751",
          4669 => x"56577474",
          4670 => x"24fac138",
          4671 => x"82cdec08",
          4672 => x"528851ff",
          4673 => x"a1ac3f74",
          4674 => x"81800a29",
          4675 => x"81800a05",
          4676 => x"70982c82",
          4677 => x"cdc83358",
          4678 => x"51557575",
          4679 => x"25de38fa",
          4680 => x"9b3982cd",
          4681 => x"c8337a05",
          4682 => x"54807434",
          4683 => x"82cdec08",
          4684 => x"528a51ff",
          4685 => x"a0fc3f82",
          4686 => x"cdc85279",
          4687 => x"51f6c93f",
          4688 => x"82b69808",
          4689 => x"81ff0654",
          4690 => x"73963882",
          4691 => x"cdc83354",
          4692 => x"73802e8f",
          4693 => x"38815373",
          4694 => x"527951f1",
          4695 => x"f33f8439",
          4696 => x"807a3480",
          4697 => x"0b82cdcc",
          4698 => x"34800b82",
          4699 => x"cdc83479",
          4700 => x"82b6980c",
          4701 => x"af3d0d04",
          4702 => x"82cdcc33",
          4703 => x"5473802e",
          4704 => x"f9ba3882",
          4705 => x"cdec0852",
          4706 => x"8851ffa0",
          4707 => x"a53f82cd",
          4708 => x"cc33ff05",
          4709 => x"547382cd",
          4710 => x"cc347381",
          4711 => x"ff0654dd",
          4712 => x"3982cdcc",
          4713 => x"3382cdc8",
          4714 => x"33555573",
          4715 => x"752ef98c",
          4716 => x"38ff1454",
          4717 => x"7382cdc8",
          4718 => x"3474982b",
          4719 => x"70982c75",
          4720 => x"81ff0656",
          4721 => x"51557474",
          4722 => x"25ad3874",
          4723 => x"1a548114",
          4724 => x"33743482",
          4725 => x"cdec0852",
          4726 => x"733351ff",
          4727 => x"9fd43f74",
          4728 => x"81800a29",
          4729 => x"81800a05",
          4730 => x"70982c82",
          4731 => x"cdc83358",
          4732 => x"51557575",
          4733 => x"24d53882",
          4734 => x"cdec0852",
          4735 => x"a051ff9f",
          4736 => x"b13f82cd",
          4737 => x"cc337098",
          4738 => x"2b70982c",
          4739 => x"82cdc833",
          4740 => x"57515657",
          4741 => x"747424f8",
          4742 => x"a33882cd",
          4743 => x"ec085288",
          4744 => x"51ff9f8e",
          4745 => x"3f748180",
          4746 => x"0a298180",
          4747 => x"0a057098",
          4748 => x"2c82cdc8",
          4749 => x"33585155",
          4750 => x"757525de",
          4751 => x"38f7fd39",
          4752 => x"82cdcc33",
          4753 => x"7081ff06",
          4754 => x"82cdc833",
          4755 => x"59565474",
          4756 => x"7727f7e8",
          4757 => x"3882cdec",
          4758 => x"08528114",
          4759 => x"547382cd",
          4760 => x"cc34741a",
          4761 => x"70335254",
          4762 => x"ff9ec73f",
          4763 => x"82cdcc33",
          4764 => x"7081ff06",
          4765 => x"82cdc833",
          4766 => x"58565475",
          4767 => x"7526d638",
          4768 => x"f7ba3982",
          4769 => x"cdcc5380",
          4770 => x"52829eec",
          4771 => x"51eef03f",
          4772 => x"800b82cd",
          4773 => x"cc34800b",
          4774 => x"82cdc834",
          4775 => x"f79e397a",
          4776 => x"b03882b5",
          4777 => x"e4085574",
          4778 => x"802ea638",
          4779 => x"7451ffa6",
          4780 => x"d43f82b6",
          4781 => x"980882cd",
          4782 => x"c83482b6",
          4783 => x"980881ff",
          4784 => x"06810553",
          4785 => x"74527951",
          4786 => x"ffa89a3f",
          4787 => x"935b81c0",
          4788 => x"397a8429",
          4789 => x"82b59805",
          4790 => x"fc110856",
          4791 => x"5474802e",
          4792 => x"a7387451",
          4793 => x"ffa69e3f",
          4794 => x"82b69808",
          4795 => x"82cdc834",
          4796 => x"82b69808",
          4797 => x"81ff0681",
          4798 => x"05537452",
          4799 => x"7951ffa7",
          4800 => x"e43fff1b",
          4801 => x"5480fa39",
          4802 => x"73085574",
          4803 => x"802ef6ac",
          4804 => x"387451ff",
          4805 => x"a5ef3f99",
          4806 => x"397a932e",
          4807 => x"098106ae",
          4808 => x"3882b598",
          4809 => x"08557480",
          4810 => x"2ea43874",
          4811 => x"51ffa5d5",
          4812 => x"3f82b698",
          4813 => x"0882cdc8",
          4814 => x"3482b698",
          4815 => x"0881ff06",
          4816 => x"81055374",
          4817 => x"527951ff",
          4818 => x"a79b3f80",
          4819 => x"c3397a84",
          4820 => x"2982b59c",
          4821 => x"05700856",
          4822 => x"5474802e",
          4823 => x"ab387451",
          4824 => x"ffa5a23f",
          4825 => x"82b69808",
          4826 => x"82cdc834",
          4827 => x"82b69808",
          4828 => x"81ff0681",
          4829 => x"05537452",
          4830 => x"7951ffa6",
          4831 => x"e83f811b",
          4832 => x"547381ff",
          4833 => x"065b8939",
          4834 => x"7482cdc8",
          4835 => x"34747a34",
          4836 => x"82cdcc53",
          4837 => x"82cdc833",
          4838 => x"527951ec",
          4839 => x"e23ff59c",
          4840 => x"3982cdcc",
          4841 => x"337081ff",
          4842 => x"0682cdc8",
          4843 => x"33595654",
          4844 => x"747727f5",
          4845 => x"873882cd",
          4846 => x"ec085281",
          4847 => x"14547382",
          4848 => x"cdcc3474",
          4849 => x"1a703352",
          4850 => x"54ff9be6",
          4851 => x"3ff4ed39",
          4852 => x"82cdcc33",
          4853 => x"5473802e",
          4854 => x"f4e23882",
          4855 => x"cdec0852",
          4856 => x"8851ff9b",
          4857 => x"cd3f82cd",
          4858 => x"cc33ff05",
          4859 => x"547382cd",
          4860 => x"cc34f4c8",
          4861 => x"39f93d0d",
          4862 => x"83bff40b",
          4863 => x"82b6900c",
          4864 => x"84800b82",
          4865 => x"b68c23a0",
          4866 => x"80538052",
          4867 => x"83bff451",
          4868 => x"ffaad33f",
          4869 => x"82b69008",
          4870 => x"54805877",
          4871 => x"74348157",
          4872 => x"76811534",
          4873 => x"82b69008",
          4874 => x"54778415",
          4875 => x"34768515",
          4876 => x"3482b690",
          4877 => x"08547786",
          4878 => x"15347687",
          4879 => x"153482b6",
          4880 => x"900882b6",
          4881 => x"8c22ff05",
          4882 => x"fe808007",
          4883 => x"7083ffff",
          4884 => x"0670882a",
          4885 => x"58515556",
          4886 => x"74881734",
          4887 => x"73891734",
          4888 => x"82b68c22",
          4889 => x"70882982",
          4890 => x"b6900805",
          4891 => x"f8115155",
          4892 => x"55778215",
          4893 => x"34768315",
          4894 => x"34893d0d",
          4895 => x"04ff3d0d",
          4896 => x"73528151",
          4897 => x"8472278f",
          4898 => x"38fb1283",
          4899 => x"2a821170",
          4900 => x"83ffff06",
          4901 => x"51515170",
          4902 => x"82b6980c",
          4903 => x"833d0d04",
          4904 => x"f93d0d02",
          4905 => x"a6052202",
          4906 => x"8405aa05",
          4907 => x"22710582",
          4908 => x"b6900871",
          4909 => x"832b7111",
          4910 => x"74832b73",
          4911 => x"11703381",
          4912 => x"12337188",
          4913 => x"2b0702a4",
          4914 => x"05ae0522",
          4915 => x"7181ffff",
          4916 => x"06077088",
          4917 => x"2a535152",
          4918 => x"59545b5b",
          4919 => x"57535455",
          4920 => x"71773470",
          4921 => x"81183482",
          4922 => x"b6900814",
          4923 => x"75882a52",
          4924 => x"54708215",
          4925 => x"34748315",
          4926 => x"3482b690",
          4927 => x"08701770",
          4928 => x"33811233",
          4929 => x"71882b07",
          4930 => x"70832b8f",
          4931 => x"fff80651",
          4932 => x"52565271",
          4933 => x"057383ff",
          4934 => x"ff067088",
          4935 => x"2a545451",
          4936 => x"71821234",
          4937 => x"7281ff06",
          4938 => x"53728312",
          4939 => x"3482b690",
          4940 => x"08165671",
          4941 => x"76347281",
          4942 => x"1734893d",
          4943 => x"0d04fb3d",
          4944 => x"0d82b690",
          4945 => x"08028405",
          4946 => x"9e052270",
          4947 => x"832b7211",
          4948 => x"86113387",
          4949 => x"1233718b",
          4950 => x"2b71832b",
          4951 => x"07585b59",
          4952 => x"52555272",
          4953 => x"05841233",
          4954 => x"85133371",
          4955 => x"882b0770",
          4956 => x"882a5456",
          4957 => x"56527084",
          4958 => x"13347385",
          4959 => x"133482b6",
          4960 => x"90087014",
          4961 => x"84113385",
          4962 => x"1233718b",
          4963 => x"2b71832b",
          4964 => x"07565957",
          4965 => x"52720586",
          4966 => x"12338713",
          4967 => x"3371882b",
          4968 => x"0770882a",
          4969 => x"54565652",
          4970 => x"70861334",
          4971 => x"73871334",
          4972 => x"82b69008",
          4973 => x"13703381",
          4974 => x"12337188",
          4975 => x"2b077081",
          4976 => x"ffff0670",
          4977 => x"882a5351",
          4978 => x"53535371",
          4979 => x"73347081",
          4980 => x"1434873d",
          4981 => x"0d04fa3d",
          4982 => x"0d02a205",
          4983 => x"2282b690",
          4984 => x"0871832b",
          4985 => x"71117033",
          4986 => x"81123371",
          4987 => x"882b0770",
          4988 => x"88291570",
          4989 => x"33811233",
          4990 => x"71982b71",
          4991 => x"902b0753",
          4992 => x"5f535552",
          4993 => x"5a565753",
          4994 => x"54718025",
          4995 => x"80f63872",
          4996 => x"51feab3f",
          4997 => x"82b69008",
          4998 => x"70167033",
          4999 => x"81123371",
          5000 => x"8b2b7183",
          5001 => x"2b077411",
          5002 => x"70338112",
          5003 => x"3371882b",
          5004 => x"0770832b",
          5005 => x"8ffff806",
          5006 => x"51525451",
          5007 => x"535a5853",
          5008 => x"72057488",
          5009 => x"2a545272",
          5010 => x"82133473",
          5011 => x"83133482",
          5012 => x"b6900870",
          5013 => x"16703381",
          5014 => x"1233718b",
          5015 => x"2b71832b",
          5016 => x"07565957",
          5017 => x"55720570",
          5018 => x"33811233",
          5019 => x"71882b07",
          5020 => x"7081ffff",
          5021 => x"0670882a",
          5022 => x"57515258",
          5023 => x"52727434",
          5024 => x"71811534",
          5025 => x"883d0d04",
          5026 => x"fb3d0d82",
          5027 => x"b6900802",
          5028 => x"84059e05",
          5029 => x"2270832b",
          5030 => x"72118211",
          5031 => x"33831233",
          5032 => x"718b2b71",
          5033 => x"832b0759",
          5034 => x"5b595256",
          5035 => x"52730571",
          5036 => x"33811333",
          5037 => x"71882b07",
          5038 => x"028c05a2",
          5039 => x"05227107",
          5040 => x"70882a53",
          5041 => x"51535353",
          5042 => x"71733470",
          5043 => x"81143482",
          5044 => x"b6900870",
          5045 => x"15703381",
          5046 => x"1233718b",
          5047 => x"2b71832b",
          5048 => x"07565957",
          5049 => x"52720582",
          5050 => x"12338313",
          5051 => x"3371882b",
          5052 => x"0770882a",
          5053 => x"54555652",
          5054 => x"70821334",
          5055 => x"72831334",
          5056 => x"82b69008",
          5057 => x"14821133",
          5058 => x"83123371",
          5059 => x"882b0782",
          5060 => x"b6980c52",
          5061 => x"54873d0d",
          5062 => x"04f73d0d",
          5063 => x"7b82b690",
          5064 => x"0831832a",
          5065 => x"7083ffff",
          5066 => x"06705357",
          5067 => x"53fda73f",
          5068 => x"82b69008",
          5069 => x"76832b71",
          5070 => x"11821133",
          5071 => x"83123371",
          5072 => x"8b2b7183",
          5073 => x"2b077511",
          5074 => x"70338112",
          5075 => x"3371982b",
          5076 => x"71902b07",
          5077 => x"53424051",
          5078 => x"535b5855",
          5079 => x"59547280",
          5080 => x"258d3882",
          5081 => x"80805275",
          5082 => x"51fe9d3f",
          5083 => x"81843984",
          5084 => x"14338515",
          5085 => x"33718b2b",
          5086 => x"71832b07",
          5087 => x"76117988",
          5088 => x"2a535155",
          5089 => x"58557686",
          5090 => x"14347581",
          5091 => x"ff065675",
          5092 => x"87143482",
          5093 => x"b6900870",
          5094 => x"19841233",
          5095 => x"85133371",
          5096 => x"882b0770",
          5097 => x"882a5457",
          5098 => x"5b565372",
          5099 => x"84163473",
          5100 => x"85163482",
          5101 => x"b6900818",
          5102 => x"53800b86",
          5103 => x"1434800b",
          5104 => x"87143482",
          5105 => x"b6900853",
          5106 => x"76841434",
          5107 => x"75851434",
          5108 => x"82b69008",
          5109 => x"18703381",
          5110 => x"12337188",
          5111 => x"2b077082",
          5112 => x"80800770",
          5113 => x"882a5351",
          5114 => x"55565474",
          5115 => x"74347281",
          5116 => x"15348b3d",
          5117 => x"0d04ff3d",
          5118 => x"0d735282",
          5119 => x"b6900884",
          5120 => x"38f7f23f",
          5121 => x"71802e86",
          5122 => x"387151fe",
          5123 => x"8c3f833d",
          5124 => x"0d04f53d",
          5125 => x"0d807e52",
          5126 => x"58f8e23f",
          5127 => x"82b69808",
          5128 => x"83ffff06",
          5129 => x"82b69008",
          5130 => x"84113385",
          5131 => x"12337188",
          5132 => x"2b07705f",
          5133 => x"5956585a",
          5134 => x"81ffff59",
          5135 => x"75782e80",
          5136 => x"cb387588",
          5137 => x"29177033",
          5138 => x"81123371",
          5139 => x"882b0770",
          5140 => x"81ffff06",
          5141 => x"79317083",
          5142 => x"ffff0670",
          5143 => x"7f275253",
          5144 => x"51565955",
          5145 => x"7779278a",
          5146 => x"3873802e",
          5147 => x"85387578",
          5148 => x"5a5b8415",
          5149 => x"33851633",
          5150 => x"71882b07",
          5151 => x"575475c2",
          5152 => x"387881ff",
          5153 => x"ff2e8538",
          5154 => x"7a795956",
          5155 => x"8076832b",
          5156 => x"82b69008",
          5157 => x"11703381",
          5158 => x"12337188",
          5159 => x"2b077081",
          5160 => x"ffff0651",
          5161 => x"525a565c",
          5162 => x"5573752e",
          5163 => x"83388155",
          5164 => x"80547978",
          5165 => x"2681cc38",
          5166 => x"74547480",
          5167 => x"2e81c438",
          5168 => x"777a2e09",
          5169 => x"81068938",
          5170 => x"7551f8f2",
          5171 => x"3f81ac39",
          5172 => x"82808053",
          5173 => x"79527551",
          5174 => x"f7c63f82",
          5175 => x"b6900870",
          5176 => x"1c861133",
          5177 => x"87123371",
          5178 => x"8b2b7183",
          5179 => x"2b07535a",
          5180 => x"5e557405",
          5181 => x"7a177083",
          5182 => x"ffff0670",
          5183 => x"882a5c59",
          5184 => x"56547884",
          5185 => x"15347681",
          5186 => x"ff065776",
          5187 => x"85153482",
          5188 => x"b6900875",
          5189 => x"832b7111",
          5190 => x"721e8611",
          5191 => x"33871233",
          5192 => x"71882b07",
          5193 => x"70882a53",
          5194 => x"5b5e535a",
          5195 => x"56547386",
          5196 => x"19347587",
          5197 => x"193482b6",
          5198 => x"9008701c",
          5199 => x"84113385",
          5200 => x"1233718b",
          5201 => x"2b71832b",
          5202 => x"07535d5a",
          5203 => x"55740554",
          5204 => x"78861534",
          5205 => x"76871534",
          5206 => x"82b69008",
          5207 => x"7016711d",
          5208 => x"84113385",
          5209 => x"12337188",
          5210 => x"2b077088",
          5211 => x"2a535a5f",
          5212 => x"52565473",
          5213 => x"84163475",
          5214 => x"85163482",
          5215 => x"b690081b",
          5216 => x"84055473",
          5217 => x"82b6980c",
          5218 => x"8d3d0d04",
          5219 => x"fe3d0d74",
          5220 => x"5282b690",
          5221 => x"088438f4",
          5222 => x"dc3f7153",
          5223 => x"71802e8b",
          5224 => x"387151fc",
          5225 => x"ed3f82b6",
          5226 => x"98085372",
          5227 => x"82b6980c",
          5228 => x"843d0d04",
          5229 => x"ee3d0d64",
          5230 => x"66405c80",
          5231 => x"70424082",
          5232 => x"b6900860",
          5233 => x"2e098106",
          5234 => x"8438f4a9",
          5235 => x"3f7b8e38",
          5236 => x"7e51ffb8",
          5237 => x"3f82b698",
          5238 => x"085483c7",
          5239 => x"397e8b38",
          5240 => x"7b51fc92",
          5241 => x"3f7e5483",
          5242 => x"ba397e51",
          5243 => x"f58f3f82",
          5244 => x"b6980883",
          5245 => x"ffff0682",
          5246 => x"b690087d",
          5247 => x"7131832a",
          5248 => x"7083ffff",
          5249 => x"0670832b",
          5250 => x"73117033",
          5251 => x"81123371",
          5252 => x"882b0770",
          5253 => x"75317083",
          5254 => x"ffff0670",
          5255 => x"8829fc05",
          5256 => x"7388291a",
          5257 => x"70338112",
          5258 => x"3371882b",
          5259 => x"0770902b",
          5260 => x"53444e53",
          5261 => x"4841525c",
          5262 => x"545b415c",
          5263 => x"565b5b73",
          5264 => x"80258f38",
          5265 => x"7681ffff",
          5266 => x"06753170",
          5267 => x"83ffff06",
          5268 => x"42548216",
          5269 => x"33831733",
          5270 => x"71882b07",
          5271 => x"7088291c",
          5272 => x"70338112",
          5273 => x"3371982b",
          5274 => x"71902b07",
          5275 => x"53474552",
          5276 => x"56547380",
          5277 => x"258b3878",
          5278 => x"75317083",
          5279 => x"ffff0641",
          5280 => x"54777b27",
          5281 => x"81fe3860",
          5282 => x"1854737b",
          5283 => x"2e098106",
          5284 => x"8f387851",
          5285 => x"f6c03f7a",
          5286 => x"83ffff06",
          5287 => x"5881e539",
          5288 => x"7f8e387a",
          5289 => x"74248938",
          5290 => x"7851f6aa",
          5291 => x"3f81a539",
          5292 => x"7f18557a",
          5293 => x"752480c8",
          5294 => x"38791d82",
          5295 => x"11338312",
          5296 => x"3371882b",
          5297 => x"07535754",
          5298 => x"f4f43f80",
          5299 => x"527851f7",
          5300 => x"b73f82b6",
          5301 => x"980883ff",
          5302 => x"ff067e54",
          5303 => x"7c537083",
          5304 => x"2b82b690",
          5305 => x"08118405",
          5306 => x"535559ff",
          5307 => x"93ad3f82",
          5308 => x"b6900814",
          5309 => x"84057583",
          5310 => x"ffff0659",
          5311 => x"5c818539",
          5312 => x"6015547a",
          5313 => x"742480d4",
          5314 => x"387851f5",
          5315 => x"c93f82b6",
          5316 => x"90081d82",
          5317 => x"11338312",
          5318 => x"3371882b",
          5319 => x"07534354",
          5320 => x"f49c3f80",
          5321 => x"527851f6",
          5322 => x"df3f82b6",
          5323 => x"980883ff",
          5324 => x"ff067e54",
          5325 => x"7c537083",
          5326 => x"2b82b690",
          5327 => x"08118405",
          5328 => x"535559ff",
          5329 => x"92d53f82",
          5330 => x"b6900814",
          5331 => x"84056062",
          5332 => x"0519555c",
          5333 => x"7383ffff",
          5334 => x"0658a939",
          5335 => x"7b7f5254",
          5336 => x"f9b03f82",
          5337 => x"b698085c",
          5338 => x"82b69808",
          5339 => x"802e9338",
          5340 => x"7d537352",
          5341 => x"82b69808",
          5342 => x"51ff96e9",
          5343 => x"3f7351f7",
          5344 => x"983f7a58",
          5345 => x"7a782799",
          5346 => x"3880537a",
          5347 => x"527851f2",
          5348 => x"8f3f7a19",
          5349 => x"832b82b6",
          5350 => x"90080584",
          5351 => x"0551f6f9",
          5352 => x"3f7b5473",
          5353 => x"82b6980c",
          5354 => x"943d0d04",
          5355 => x"fc3d0d77",
          5356 => x"77297052",
          5357 => x"54fbd53f",
          5358 => x"82b69808",
          5359 => x"5582b698",
          5360 => x"08802e8e",
          5361 => x"38735380",
          5362 => x"5282b698",
          5363 => x"0851ff9b",
          5364 => x"953f7482",
          5365 => x"b6980c86",
          5366 => x"3d0d04ff",
          5367 => x"3d0d028f",
          5368 => x"05335181",
          5369 => x"52707226",
          5370 => x"873882b6",
          5371 => x"94113352",
          5372 => x"7182b698",
          5373 => x"0c833d0d",
          5374 => x"04fc3d0d",
          5375 => x"029b0533",
          5376 => x"0284059f",
          5377 => x"05335653",
          5378 => x"83517281",
          5379 => x"2680e038",
          5380 => x"72842b87",
          5381 => x"c0928c11",
          5382 => x"53518854",
          5383 => x"74802e84",
          5384 => x"38818854",
          5385 => x"73720c87",
          5386 => x"c0928c11",
          5387 => x"5181710c",
          5388 => x"850b87c0",
          5389 => x"988c0c70",
          5390 => x"52710870",
          5391 => x"82065151",
          5392 => x"70802e8a",
          5393 => x"3887c098",
          5394 => x"8c085170",
          5395 => x"ec387108",
          5396 => x"fc808006",
          5397 => x"52719238",
          5398 => x"87c0988c",
          5399 => x"08517080",
          5400 => x"2e873871",
          5401 => x"82b69414",
          5402 => x"3482b694",
          5403 => x"13335170",
          5404 => x"82b6980c",
          5405 => x"863d0d04",
          5406 => x"f33d0d60",
          5407 => x"6264028c",
          5408 => x"05bf0533",
          5409 => x"5740585b",
          5410 => x"8374525a",
          5411 => x"fecd3f82",
          5412 => x"b6980881",
          5413 => x"067a5452",
          5414 => x"7181be38",
          5415 => x"71727584",
          5416 => x"2b87c092",
          5417 => x"801187c0",
          5418 => x"928c1287",
          5419 => x"c0928413",
          5420 => x"415a4057",
          5421 => x"5a58850b",
          5422 => x"87c0988c",
          5423 => x"0c767d0c",
          5424 => x"84760c75",
          5425 => x"0870852a",
          5426 => x"70810651",
          5427 => x"53547180",
          5428 => x"2e8e387b",
          5429 => x"0852717b",
          5430 => x"7081055d",
          5431 => x"34811959",
          5432 => x"8074a206",
          5433 => x"53537173",
          5434 => x"2e833881",
          5435 => x"537883ff",
          5436 => x"268f3872",
          5437 => x"802e8a38",
          5438 => x"87c0988c",
          5439 => x"085271c3",
          5440 => x"3887c098",
          5441 => x"8c085271",
          5442 => x"802e8738",
          5443 => x"7884802e",
          5444 => x"99388176",
          5445 => x"0c87c092",
          5446 => x"8c155372",
          5447 => x"08708206",
          5448 => x"515271f7",
          5449 => x"38ff1a5a",
          5450 => x"8d398480",
          5451 => x"17811970",
          5452 => x"81ff065a",
          5453 => x"53577980",
          5454 => x"2e903873",
          5455 => x"fc808006",
          5456 => x"52718738",
          5457 => x"7d7826fe",
          5458 => x"ed3873fc",
          5459 => x"80800652",
          5460 => x"71802e83",
          5461 => x"38815271",
          5462 => x"537282b6",
          5463 => x"980c8f3d",
          5464 => x"0d04f33d",
          5465 => x"0d606264",
          5466 => x"028c05bf",
          5467 => x"05335740",
          5468 => x"585b8359",
          5469 => x"80745258",
          5470 => x"fce13f82",
          5471 => x"b6980881",
          5472 => x"06795452",
          5473 => x"71782e09",
          5474 => x"810681b1",
          5475 => x"38777484",
          5476 => x"2b87c092",
          5477 => x"801187c0",
          5478 => x"928c1287",
          5479 => x"c0928413",
          5480 => x"40595f56",
          5481 => x"5a850b87",
          5482 => x"c0988c0c",
          5483 => x"767d0c82",
          5484 => x"760c8058",
          5485 => x"75087084",
          5486 => x"2a708106",
          5487 => x"51535471",
          5488 => x"802e8c38",
          5489 => x"7a708105",
          5490 => x"5c337c0c",
          5491 => x"81185873",
          5492 => x"812a7081",
          5493 => x"06515271",
          5494 => x"802e8a38",
          5495 => x"87c0988c",
          5496 => x"085271d0",
          5497 => x"3887c098",
          5498 => x"8c085271",
          5499 => x"802e8738",
          5500 => x"7784802e",
          5501 => x"99388176",
          5502 => x"0c87c092",
          5503 => x"8c155372",
          5504 => x"08708206",
          5505 => x"515271f7",
          5506 => x"38ff1959",
          5507 => x"8d39811a",
          5508 => x"7081ff06",
          5509 => x"84801959",
          5510 => x"5b527880",
          5511 => x"2e903873",
          5512 => x"fc808006",
          5513 => x"52718738",
          5514 => x"7d7a26fe",
          5515 => x"f83873fc",
          5516 => x"80800652",
          5517 => x"71802e83",
          5518 => x"38815271",
          5519 => x"537282b6",
          5520 => x"980c8f3d",
          5521 => x"0d04fa3d",
          5522 => x"0d7a0284",
          5523 => x"05a30533",
          5524 => x"028805a7",
          5525 => x"05337154",
          5526 => x"545657fa",
          5527 => x"fe3f82b6",
          5528 => x"98088106",
          5529 => x"53835472",
          5530 => x"80fe3885",
          5531 => x"0b87c098",
          5532 => x"8c0c8156",
          5533 => x"71762e80",
          5534 => x"dc387176",
          5535 => x"24933874",
          5536 => x"842b87c0",
          5537 => x"928c1154",
          5538 => x"5471802e",
          5539 => x"8d3880d4",
          5540 => x"3971832e",
          5541 => x"80c63880",
          5542 => x"cb397208",
          5543 => x"70812a70",
          5544 => x"81065151",
          5545 => x"5271802e",
          5546 => x"8a3887c0",
          5547 => x"988c0852",
          5548 => x"71e83887",
          5549 => x"c0988c08",
          5550 => x"52719638",
          5551 => x"81730c87",
          5552 => x"c0928c14",
          5553 => x"53720870",
          5554 => x"82065152",
          5555 => x"71f73896",
          5556 => x"39805692",
          5557 => x"3988800a",
          5558 => x"770c8539",
          5559 => x"8180770c",
          5560 => x"72568339",
          5561 => x"84567554",
          5562 => x"7382b698",
          5563 => x"0c883d0d",
          5564 => x"04fe3d0d",
          5565 => x"74811133",
          5566 => x"71337188",
          5567 => x"2b0782b6",
          5568 => x"980c5351",
          5569 => x"843d0d04",
          5570 => x"fd3d0d75",
          5571 => x"83113382",
          5572 => x"12337190",
          5573 => x"2b71882b",
          5574 => x"07811433",
          5575 => x"70720788",
          5576 => x"2b753371",
          5577 => x"0782b698",
          5578 => x"0c525354",
          5579 => x"56545285",
          5580 => x"3d0d04ff",
          5581 => x"3d0d7302",
          5582 => x"84059205",
          5583 => x"22525270",
          5584 => x"72708105",
          5585 => x"54347088",
          5586 => x"2a517072",
          5587 => x"34833d0d",
          5588 => x"04ff3d0d",
          5589 => x"73755252",
          5590 => x"70727081",
          5591 => x"05543470",
          5592 => x"882a5170",
          5593 => x"72708105",
          5594 => x"54347088",
          5595 => x"2a517072",
          5596 => x"70810554",
          5597 => x"3470882a",
          5598 => x"51707234",
          5599 => x"833d0d04",
          5600 => x"fe3d0d76",
          5601 => x"75775454",
          5602 => x"5170802e",
          5603 => x"92387170",
          5604 => x"81055333",
          5605 => x"73708105",
          5606 => x"5534ff11",
          5607 => x"51eb3984",
          5608 => x"3d0d04fe",
          5609 => x"3d0d7577",
          5610 => x"76545253",
          5611 => x"72727081",
          5612 => x"055434ff",
          5613 => x"115170f4",
          5614 => x"38843d0d",
          5615 => x"04fc3d0d",
          5616 => x"78777956",
          5617 => x"56537470",
          5618 => x"81055633",
          5619 => x"74708105",
          5620 => x"56337171",
          5621 => x"31ff1656",
          5622 => x"52525272",
          5623 => x"802e8638",
          5624 => x"71802ee2",
          5625 => x"387182b6",
          5626 => x"980c863d",
          5627 => x"0d04fe3d",
          5628 => x"0d747654",
          5629 => x"51893971",
          5630 => x"732e8a38",
          5631 => x"81115170",
          5632 => x"335271f3",
          5633 => x"38703382",
          5634 => x"b6980c84",
          5635 => x"3d0d0480",
          5636 => x"0b82b698",
          5637 => x"0c04800b",
          5638 => x"82b6980c",
          5639 => x"04f73d0d",
          5640 => x"7b56800b",
          5641 => x"83173356",
          5642 => x"5a747a2e",
          5643 => x"80d63881",
          5644 => x"54b01608",
          5645 => x"53b41670",
          5646 => x"53811733",
          5647 => x"5259faa2",
          5648 => x"3f82b698",
          5649 => x"087a2e09",
          5650 => x"8106b738",
          5651 => x"82b69808",
          5652 => x"831734b0",
          5653 => x"160870a4",
          5654 => x"1808319c",
          5655 => x"18085956",
          5656 => x"58747727",
          5657 => x"9f388216",
          5658 => x"33557482",
          5659 => x"2e098106",
          5660 => x"93388154",
          5661 => x"76185378",
          5662 => x"52811633",
          5663 => x"51f9e33f",
          5664 => x"8339815a",
          5665 => x"7982b698",
          5666 => x"0c8b3d0d",
          5667 => x"04fa3d0d",
          5668 => x"787a5656",
          5669 => x"805774b0",
          5670 => x"17082eaf",
          5671 => x"387551fe",
          5672 => x"fc3f82b6",
          5673 => x"98085782",
          5674 => x"b698089f",
          5675 => x"38815474",
          5676 => x"53b41652",
          5677 => x"81163351",
          5678 => x"f7be3f82",
          5679 => x"b6980880",
          5680 => x"2e8538ff",
          5681 => x"55815774",
          5682 => x"b0170c76",
          5683 => x"82b6980c",
          5684 => x"883d0d04",
          5685 => x"f83d0d7a",
          5686 => x"705257fe",
          5687 => x"c03f82b6",
          5688 => x"98085882",
          5689 => x"b6980881",
          5690 => x"91387633",
          5691 => x"5574832e",
          5692 => x"09810680",
          5693 => x"f0388417",
          5694 => x"33597881",
          5695 => x"2e098106",
          5696 => x"80e33884",
          5697 => x"805382b6",
          5698 => x"980852b4",
          5699 => x"17705256",
          5700 => x"fd913f82",
          5701 => x"d4d55284",
          5702 => x"b21751fc",
          5703 => x"963f848b",
          5704 => x"85a4d252",
          5705 => x"7551fca9",
          5706 => x"3f868a85",
          5707 => x"e4f25284",
          5708 => x"981751fc",
          5709 => x"9c3f9017",
          5710 => x"0852849c",
          5711 => x"1751fc91",
          5712 => x"3f8c1708",
          5713 => x"5284a017",
          5714 => x"51fc863f",
          5715 => x"a0170881",
          5716 => x"0570b019",
          5717 => x"0c795553",
          5718 => x"75528117",
          5719 => x"3351f882",
          5720 => x"3f778418",
          5721 => x"34805380",
          5722 => x"52811733",
          5723 => x"51f9d73f",
          5724 => x"82b69808",
          5725 => x"802e8338",
          5726 => x"81587782",
          5727 => x"b6980c8a",
          5728 => x"3d0d04fb",
          5729 => x"3d0d77fe",
          5730 => x"1a981208",
          5731 => x"fe055556",
          5732 => x"54805674",
          5733 => x"73278d38",
          5734 => x"8a142275",
          5735 => x"7129ac16",
          5736 => x"08055753",
          5737 => x"7582b698",
          5738 => x"0c873d0d",
          5739 => x"04f93d0d",
          5740 => x"7a7a7008",
          5741 => x"56545781",
          5742 => x"772781df",
          5743 => x"38769815",
          5744 => x"082781d7",
          5745 => x"38ff7433",
          5746 => x"54587282",
          5747 => x"2e80f538",
          5748 => x"72822489",
          5749 => x"3872812e",
          5750 => x"8d3881bf",
          5751 => x"3972832e",
          5752 => x"818e3881",
          5753 => x"b6397681",
          5754 => x"2a177089",
          5755 => x"2aa41608",
          5756 => x"05537452",
          5757 => x"55fd963f",
          5758 => x"82b69808",
          5759 => x"819f3874",
          5760 => x"83ff0614",
          5761 => x"b4113381",
          5762 => x"1770892a",
          5763 => x"a4180805",
          5764 => x"55765457",
          5765 => x"5753fcf5",
          5766 => x"3f82b698",
          5767 => x"0880fe38",
          5768 => x"7483ff06",
          5769 => x"14b41133",
          5770 => x"70882b78",
          5771 => x"07798106",
          5772 => x"71842a5c",
          5773 => x"52585153",
          5774 => x"7280e238",
          5775 => x"759fff06",
          5776 => x"5880da39",
          5777 => x"76882aa4",
          5778 => x"15080552",
          5779 => x"7351fcbd",
          5780 => x"3f82b698",
          5781 => x"0880c638",
          5782 => x"761083fe",
          5783 => x"067405b4",
          5784 => x"0551f98d",
          5785 => x"3f82b698",
          5786 => x"0883ffff",
          5787 => x"0658ae39",
          5788 => x"76872aa4",
          5789 => x"15080552",
          5790 => x"7351fc91",
          5791 => x"3f82b698",
          5792 => x"089b3876",
          5793 => x"822b83fc",
          5794 => x"067405b4",
          5795 => x"0551f8f8",
          5796 => x"3f82b698",
          5797 => x"08f00a06",
          5798 => x"58833981",
          5799 => x"587782b6",
          5800 => x"980c893d",
          5801 => x"0d04f83d",
          5802 => x"0d7a7c7e",
          5803 => x"5a585682",
          5804 => x"59817727",
          5805 => x"829e3876",
          5806 => x"98170827",
          5807 => x"82963875",
          5808 => x"33537279",
          5809 => x"2e819d38",
          5810 => x"72792489",
          5811 => x"3872812e",
          5812 => x"8d388280",
          5813 => x"3972832e",
          5814 => x"81b83881",
          5815 => x"f7397681",
          5816 => x"2a177089",
          5817 => x"2aa41808",
          5818 => x"05537652",
          5819 => x"55fb9e3f",
          5820 => x"82b69808",
          5821 => x"5982b698",
          5822 => x"0881d938",
          5823 => x"7483ff06",
          5824 => x"16b40581",
          5825 => x"16788106",
          5826 => x"59565477",
          5827 => x"5376802e",
          5828 => x"8f387784",
          5829 => x"2b9ff006",
          5830 => x"74338f06",
          5831 => x"71075153",
          5832 => x"72743481",
          5833 => x"0b831734",
          5834 => x"74892aa4",
          5835 => x"17080552",
          5836 => x"7551fad9",
          5837 => x"3f82b698",
          5838 => x"085982b6",
          5839 => x"98088194",
          5840 => x"387483ff",
          5841 => x"0616b405",
          5842 => x"78842a54",
          5843 => x"54768f38",
          5844 => x"77882a74",
          5845 => x"3381f006",
          5846 => x"718f0607",
          5847 => x"51537274",
          5848 => x"3480ec39",
          5849 => x"76882aa4",
          5850 => x"17080552",
          5851 => x"7551fa9d",
          5852 => x"3f82b698",
          5853 => x"085982b6",
          5854 => x"980880d8",
          5855 => x"387783ff",
          5856 => x"ff065276",
          5857 => x"1083fe06",
          5858 => x"7605b405",
          5859 => x"51f7a43f",
          5860 => x"be397687",
          5861 => x"2aa41708",
          5862 => x"05527551",
          5863 => x"f9ef3f82",
          5864 => x"b6980859",
          5865 => x"82b69808",
          5866 => x"ab3877f0",
          5867 => x"0a067782",
          5868 => x"2b83fc06",
          5869 => x"7018b405",
          5870 => x"70545154",
          5871 => x"54f6c93f",
          5872 => x"82b69808",
          5873 => x"8f0a0674",
          5874 => x"07527251",
          5875 => x"f7833f81",
          5876 => x"0b831734",
          5877 => x"7882b698",
          5878 => x"0c8a3d0d",
          5879 => x"04f83d0d",
          5880 => x"7a7c7e72",
          5881 => x"08595656",
          5882 => x"59817527",
          5883 => x"a4387498",
          5884 => x"1708279d",
          5885 => x"3873802e",
          5886 => x"aa38ff53",
          5887 => x"73527551",
          5888 => x"fda43f82",
          5889 => x"b6980854",
          5890 => x"82b69808",
          5891 => x"80f23893",
          5892 => x"39825480",
          5893 => x"eb398154",
          5894 => x"80e63982",
          5895 => x"b6980854",
          5896 => x"80de3974",
          5897 => x"527851fb",
          5898 => x"843f82b6",
          5899 => x"98085882",
          5900 => x"b6980880",
          5901 => x"2e80c738",
          5902 => x"82b69808",
          5903 => x"812ed238",
          5904 => x"82b69808",
          5905 => x"ff2ecf38",
          5906 => x"80537452",
          5907 => x"7551fcd6",
          5908 => x"3f82b698",
          5909 => x"08c53898",
          5910 => x"1608fe11",
          5911 => x"90180857",
          5912 => x"55577474",
          5913 => x"27903881",
          5914 => x"1590170c",
          5915 => x"84163381",
          5916 => x"07547384",
          5917 => x"17347755",
          5918 => x"767826ff",
          5919 => x"a6388054",
          5920 => x"7382b698",
          5921 => x"0c8a3d0d",
          5922 => x"04f63d0d",
          5923 => x"7c7e7108",
          5924 => x"595b5b79",
          5925 => x"95388c17",
          5926 => x"08587780",
          5927 => x"2e883898",
          5928 => x"17087826",
          5929 => x"b2388158",
          5930 => x"ae397952",
          5931 => x"7a51f9fd",
          5932 => x"3f815574",
          5933 => x"82b69808",
          5934 => x"2782e038",
          5935 => x"82b69808",
          5936 => x"5582b698",
          5937 => x"08ff2e82",
          5938 => x"d2389817",
          5939 => x"0882b698",
          5940 => x"082682c7",
          5941 => x"38795890",
          5942 => x"17087056",
          5943 => x"5473802e",
          5944 => x"82b93877",
          5945 => x"7a2e0981",
          5946 => x"0680e238",
          5947 => x"811a5698",
          5948 => x"17087626",
          5949 => x"83388256",
          5950 => x"75527a51",
          5951 => x"f9af3f80",
          5952 => x"5982b698",
          5953 => x"08812e09",
          5954 => x"81068638",
          5955 => x"82b69808",
          5956 => x"5982b698",
          5957 => x"08097030",
          5958 => x"70720780",
          5959 => x"25707c07",
          5960 => x"82b69808",
          5961 => x"54515155",
          5962 => x"557381ef",
          5963 => x"3882b698",
          5964 => x"08802e95",
          5965 => x"388c1708",
          5966 => x"54817427",
          5967 => x"90387398",
          5968 => x"18082789",
          5969 => x"38735885",
          5970 => x"397580db",
          5971 => x"38775681",
          5972 => x"16569817",
          5973 => x"08762689",
          5974 => x"38825675",
          5975 => x"782681ac",
          5976 => x"3875527a",
          5977 => x"51f8c63f",
          5978 => x"82b69808",
          5979 => x"802eb838",
          5980 => x"805982b6",
          5981 => x"9808812e",
          5982 => x"09810686",
          5983 => x"3882b698",
          5984 => x"085982b6",
          5985 => x"98080970",
          5986 => x"30707207",
          5987 => x"8025707c",
          5988 => x"07515155",
          5989 => x"557380f8",
          5990 => x"3875782e",
          5991 => x"098106ff",
          5992 => x"ae387355",
          5993 => x"80f539ff",
          5994 => x"53755276",
          5995 => x"51f9f73f",
          5996 => x"82b69808",
          5997 => x"82b69808",
          5998 => x"307082b6",
          5999 => x"98080780",
          6000 => x"25515555",
          6001 => x"79802e94",
          6002 => x"3873802e",
          6003 => x"8f387553",
          6004 => x"79527651",
          6005 => x"f9d03f82",
          6006 => x"b6980855",
          6007 => x"74a53875",
          6008 => x"8c180c98",
          6009 => x"1708fe05",
          6010 => x"90180856",
          6011 => x"54747426",
          6012 => x"8638ff15",
          6013 => x"90180c84",
          6014 => x"17338107",
          6015 => x"54738418",
          6016 => x"349739ff",
          6017 => x"5674812e",
          6018 => x"90388c39",
          6019 => x"80558c39",
          6020 => x"82b69808",
          6021 => x"55853981",
          6022 => x"56755574",
          6023 => x"82b6980c",
          6024 => x"8c3d0d04",
          6025 => x"f83d0d7a",
          6026 => x"705255f3",
          6027 => x"f03f82b6",
          6028 => x"98085881",
          6029 => x"5682b698",
          6030 => x"0880d838",
          6031 => x"7b527451",
          6032 => x"f6c13f82",
          6033 => x"b6980882",
          6034 => x"b69808b0",
          6035 => x"170c5984",
          6036 => x"80537752",
          6037 => x"b4157052",
          6038 => x"57f2c83f",
          6039 => x"77568439",
          6040 => x"8116568a",
          6041 => x"15225875",
          6042 => x"78279738",
          6043 => x"81547519",
          6044 => x"53765281",
          6045 => x"153351ed",
          6046 => x"e93f82b6",
          6047 => x"9808802e",
          6048 => x"df388a15",
          6049 => x"22763270",
          6050 => x"30707207",
          6051 => x"709f2a53",
          6052 => x"51565675",
          6053 => x"82b6980c",
          6054 => x"8a3d0d04",
          6055 => x"f83d0d7a",
          6056 => x"7c710858",
          6057 => x"565774f0",
          6058 => x"800a2680",
          6059 => x"f138749f",
          6060 => x"06537280",
          6061 => x"e9387490",
          6062 => x"180c8817",
          6063 => x"085473aa",
          6064 => x"38753353",
          6065 => x"82732788",
          6066 => x"38a81608",
          6067 => x"54739b38",
          6068 => x"74852a53",
          6069 => x"820b8817",
          6070 => x"225a5872",
          6071 => x"792780fe",
          6072 => x"38a81608",
          6073 => x"98180c80",
          6074 => x"cd398a16",
          6075 => x"2270892b",
          6076 => x"54587275",
          6077 => x"26b23873",
          6078 => x"527651f5",
          6079 => x"b03f82b6",
          6080 => x"98085482",
          6081 => x"b69808ff",
          6082 => x"2ebd3881",
          6083 => x"0b82b698",
          6084 => x"08278b38",
          6085 => x"98160882",
          6086 => x"b6980826",
          6087 => x"85388258",
          6088 => x"bd397473",
          6089 => x"3155cb39",
          6090 => x"73527551",
          6091 => x"f4d53f82",
          6092 => x"b6980898",
          6093 => x"180c7394",
          6094 => x"180c9817",
          6095 => x"08538258",
          6096 => x"72802e9a",
          6097 => x"38853981",
          6098 => x"58943974",
          6099 => x"892a1398",
          6100 => x"180c7483",
          6101 => x"ff0616b4",
          6102 => x"059c180c",
          6103 => x"80587782",
          6104 => x"b6980c8a",
          6105 => x"3d0d04f8",
          6106 => x"3d0d7a70",
          6107 => x"08901208",
          6108 => x"a0055957",
          6109 => x"54f0800a",
          6110 => x"77278638",
          6111 => x"800b9815",
          6112 => x"0c981408",
          6113 => x"53845572",
          6114 => x"802e81cb",
          6115 => x"387683ff",
          6116 => x"06587781",
          6117 => x"b5388113",
          6118 => x"98150c94",
          6119 => x"14085574",
          6120 => x"92387685",
          6121 => x"2a881722",
          6122 => x"56537473",
          6123 => x"26819b38",
          6124 => x"80c0398a",
          6125 => x"1622ff05",
          6126 => x"77892a06",
          6127 => x"5372818a",
          6128 => x"38745273",
          6129 => x"51f3e63f",
          6130 => x"82b69808",
          6131 => x"53825581",
          6132 => x"0b82b698",
          6133 => x"082780ff",
          6134 => x"38815582",
          6135 => x"b69808ff",
          6136 => x"2e80f438",
          6137 => x"98160882",
          6138 => x"b6980826",
          6139 => x"80ca387b",
          6140 => x"8a387798",
          6141 => x"150c8455",
          6142 => x"80dd3994",
          6143 => x"14085273",
          6144 => x"51f9863f",
          6145 => x"82b69808",
          6146 => x"53875582",
          6147 => x"b6980880",
          6148 => x"2e80c438",
          6149 => x"825582b6",
          6150 => x"9808812e",
          6151 => x"ba388155",
          6152 => x"82b69808",
          6153 => x"ff2eb038",
          6154 => x"82b69808",
          6155 => x"527551fb",
          6156 => x"f33f82b6",
          6157 => x"9808a038",
          6158 => x"7294150c",
          6159 => x"72527551",
          6160 => x"f2c13f82",
          6161 => x"b6980898",
          6162 => x"150c7690",
          6163 => x"150c7716",
          6164 => x"b4059c15",
          6165 => x"0c805574",
          6166 => x"82b6980c",
          6167 => x"8a3d0d04",
          6168 => x"f73d0d7b",
          6169 => x"7d71085b",
          6170 => x"5b578052",
          6171 => x"7651fcac",
          6172 => x"3f82b698",
          6173 => x"085482b6",
          6174 => x"980880ec",
          6175 => x"3882b698",
          6176 => x"08569817",
          6177 => x"08527851",
          6178 => x"f0833f82",
          6179 => x"b6980854",
          6180 => x"82b69808",
          6181 => x"80d23882",
          6182 => x"b698089c",
          6183 => x"18087033",
          6184 => x"51545872",
          6185 => x"81e52e09",
          6186 => x"81068338",
          6187 => x"815882b6",
          6188 => x"98085572",
          6189 => x"83388155",
          6190 => x"77750753",
          6191 => x"72802e8e",
          6192 => x"38811656",
          6193 => x"757a2e09",
          6194 => x"81068838",
          6195 => x"a53982b6",
          6196 => x"98085681",
          6197 => x"527651fd",
          6198 => x"8e3f82b6",
          6199 => x"98085482",
          6200 => x"b6980880",
          6201 => x"2eff9b38",
          6202 => x"73842e09",
          6203 => x"81068338",
          6204 => x"87547382",
          6205 => x"b6980c8b",
          6206 => x"3d0d04fd",
          6207 => x"3d0d769a",
          6208 => x"115254eb",
          6209 => x"ec3f82b6",
          6210 => x"980883ff",
          6211 => x"ff067670",
          6212 => x"33515353",
          6213 => x"71832e09",
          6214 => x"81069038",
          6215 => x"941451eb",
          6216 => x"d03f82b6",
          6217 => x"9808902b",
          6218 => x"73075372",
          6219 => x"82b6980c",
          6220 => x"853d0d04",
          6221 => x"fc3d0d77",
          6222 => x"797083ff",
          6223 => x"ff06549a",
          6224 => x"12535555",
          6225 => x"ebed3f76",
          6226 => x"70335153",
          6227 => x"72832e09",
          6228 => x"81068b38",
          6229 => x"73902a52",
          6230 => x"941551eb",
          6231 => x"d63f863d",
          6232 => x"0d04f73d",
          6233 => x"0d7b7d5b",
          6234 => x"55847508",
          6235 => x"5a589815",
          6236 => x"08802e81",
          6237 => x"8a389815",
          6238 => x"08527851",
          6239 => x"ee8f3f82",
          6240 => x"b6980858",
          6241 => x"82b69808",
          6242 => x"80f5389c",
          6243 => x"15087033",
          6244 => x"55537386",
          6245 => x"38845880",
          6246 => x"e6398b13",
          6247 => x"3370bf06",
          6248 => x"7081ff06",
          6249 => x"58515372",
          6250 => x"86163482",
          6251 => x"b6980853",
          6252 => x"7381e52e",
          6253 => x"83388153",
          6254 => x"73ae2ea9",
          6255 => x"38817074",
          6256 => x"06545772",
          6257 => x"802e9e38",
          6258 => x"758f2e99",
          6259 => x"3882b698",
          6260 => x"0876df06",
          6261 => x"54547288",
          6262 => x"2e098106",
          6263 => x"83387654",
          6264 => x"737a2ea0",
          6265 => x"38805274",
          6266 => x"51fafc3f",
          6267 => x"82b69808",
          6268 => x"5882b698",
          6269 => x"08893898",
          6270 => x"1508fefa",
          6271 => x"38863980",
          6272 => x"0b98160c",
          6273 => x"7782b698",
          6274 => x"0c8b3d0d",
          6275 => x"04fb3d0d",
          6276 => x"77700857",
          6277 => x"54815273",
          6278 => x"51fcc53f",
          6279 => x"82b69808",
          6280 => x"5582b698",
          6281 => x"08b43898",
          6282 => x"14085275",
          6283 => x"51ecde3f",
          6284 => x"82b69808",
          6285 => x"5582b698",
          6286 => x"08a038a0",
          6287 => x"5382b698",
          6288 => x"08529c14",
          6289 => x"0851eadb",
          6290 => x"3f8b53a0",
          6291 => x"14529c14",
          6292 => x"0851eaac",
          6293 => x"3f810b83",
          6294 => x"17347482",
          6295 => x"b6980c87",
          6296 => x"3d0d04fd",
          6297 => x"3d0d7570",
          6298 => x"08981208",
          6299 => x"54705355",
          6300 => x"53ec9a3f",
          6301 => x"82b69808",
          6302 => x"8d389c13",
          6303 => x"0853e573",
          6304 => x"34810b83",
          6305 => x"1534853d",
          6306 => x"0d04fa3d",
          6307 => x"0d787a57",
          6308 => x"57800b89",
          6309 => x"17349817",
          6310 => x"08802e81",
          6311 => x"82388070",
          6312 => x"89185555",
          6313 => x"559c1708",
          6314 => x"14703381",
          6315 => x"16565152",
          6316 => x"71a02ea8",
          6317 => x"3871852e",
          6318 => x"09810684",
          6319 => x"3881e552",
          6320 => x"73892e09",
          6321 => x"81068b38",
          6322 => x"ae737081",
          6323 => x"05553481",
          6324 => x"15557173",
          6325 => x"70810555",
          6326 => x"34811555",
          6327 => x"8a7427c5",
          6328 => x"38751588",
          6329 => x"0552800b",
          6330 => x"8113349c",
          6331 => x"1708528b",
          6332 => x"12338817",
          6333 => x"349c1708",
          6334 => x"9c115252",
          6335 => x"e88a3f82",
          6336 => x"b6980876",
          6337 => x"0c961251",
          6338 => x"e7e73f82",
          6339 => x"b6980886",
          6340 => x"17239812",
          6341 => x"51e7da3f",
          6342 => x"82b69808",
          6343 => x"84172388",
          6344 => x"3d0d04f3",
          6345 => x"3d0d7f70",
          6346 => x"085e5b80",
          6347 => x"61703351",
          6348 => x"555573af",
          6349 => x"2e833881",
          6350 => x"557380dc",
          6351 => x"2e913874",
          6352 => x"802e8c38",
          6353 => x"941d0888",
          6354 => x"1c0caa39",
          6355 => x"81154180",
          6356 => x"61703356",
          6357 => x"565673af",
          6358 => x"2e098106",
          6359 => x"83388156",
          6360 => x"7380dc32",
          6361 => x"70307080",
          6362 => x"25780751",
          6363 => x"515473dc",
          6364 => x"3873881c",
          6365 => x"0c607033",
          6366 => x"5154739f",
          6367 => x"269638ff",
          6368 => x"800bab1c",
          6369 => x"3480527a",
          6370 => x"51f6913f",
          6371 => x"82b69808",
          6372 => x"55859839",
          6373 => x"913d61a0",
          6374 => x"1d5c5a5e",
          6375 => x"8b53a052",
          6376 => x"7951e7ff",
          6377 => x"3f807059",
          6378 => x"57887933",
          6379 => x"555c73ae",
          6380 => x"2e098106",
          6381 => x"80d43878",
          6382 => x"18703381",
          6383 => x"1a71ae32",
          6384 => x"7030709f",
          6385 => x"2a738226",
          6386 => x"07515153",
          6387 => x"5a575473",
          6388 => x"8c387917",
          6389 => x"54757434",
          6390 => x"811757db",
          6391 => x"3975af32",
          6392 => x"7030709f",
          6393 => x"2a515154",
          6394 => x"7580dc2e",
          6395 => x"8c387380",
          6396 => x"2e873875",
          6397 => x"a02682bd",
          6398 => x"3877197e",
          6399 => x"0ca454a0",
          6400 => x"762782bd",
          6401 => x"38a05482",
          6402 => x"b8397818",
          6403 => x"7033811a",
          6404 => x"5a5754a0",
          6405 => x"762781fc",
          6406 => x"3875af32",
          6407 => x"70307780",
          6408 => x"dc327030",
          6409 => x"72802571",
          6410 => x"80250751",
          6411 => x"51565155",
          6412 => x"73802eac",
          6413 => x"38843981",
          6414 => x"18588078",
          6415 => x"1a703351",
          6416 => x"555573af",
          6417 => x"2e098106",
          6418 => x"83388155",
          6419 => x"7380dc32",
          6420 => x"70307080",
          6421 => x"25770751",
          6422 => x"515473db",
          6423 => x"3881b539",
          6424 => x"75ae2e09",
          6425 => x"81068338",
          6426 => x"8154767c",
          6427 => x"27740754",
          6428 => x"73802ea2",
          6429 => x"387b8b32",
          6430 => x"703077ae",
          6431 => x"32703072",
          6432 => x"8025719f",
          6433 => x"2a075351",
          6434 => x"56515574",
          6435 => x"81a73888",
          6436 => x"578b5cfe",
          6437 => x"f5397598",
          6438 => x"2b547380",
          6439 => x"258c3875",
          6440 => x"80ff0682",
          6441 => x"afe01133",
          6442 => x"57547551",
          6443 => x"e6e13f82",
          6444 => x"b6980880",
          6445 => x"2eb23878",
          6446 => x"18703381",
          6447 => x"1a71545a",
          6448 => x"5654e6d2",
          6449 => x"3f82b698",
          6450 => x"08802e80",
          6451 => x"e838ff1c",
          6452 => x"54767427",
          6453 => x"80df3879",
          6454 => x"17547574",
          6455 => x"3481177a",
          6456 => x"11555774",
          6457 => x"7434a739",
          6458 => x"755282af",
          6459 => x"8051e5fe",
          6460 => x"3f82b698",
          6461 => x"08bf38ff",
          6462 => x"9f165473",
          6463 => x"99268938",
          6464 => x"e0167081",
          6465 => x"ff065754",
          6466 => x"79175475",
          6467 => x"74348117",
          6468 => x"57fdf739",
          6469 => x"77197e0c",
          6470 => x"76802e99",
          6471 => x"38793354",
          6472 => x"7381e52e",
          6473 => x"09810684",
          6474 => x"38857a34",
          6475 => x"8454a076",
          6476 => x"278f388b",
          6477 => x"39865581",
          6478 => x"f2398456",
          6479 => x"80f33980",
          6480 => x"54738b1b",
          6481 => x"34807b08",
          6482 => x"58527a51",
          6483 => x"f2ce3f82",
          6484 => x"b6980856",
          6485 => x"82b69808",
          6486 => x"80d73898",
          6487 => x"1b085276",
          6488 => x"51e6aa3f",
          6489 => x"82b69808",
          6490 => x"5682b698",
          6491 => x"0880c238",
          6492 => x"9c1b0870",
          6493 => x"33555573",
          6494 => x"802effbe",
          6495 => x"388b1533",
          6496 => x"bf065473",
          6497 => x"861c348b",
          6498 => x"15337083",
          6499 => x"2a708106",
          6500 => x"51555873",
          6501 => x"92388b53",
          6502 => x"79527451",
          6503 => x"e49f3f82",
          6504 => x"b6980880",
          6505 => x"2e8b3875",
          6506 => x"527a51f3",
          6507 => x"ba3fff9f",
          6508 => x"3975ab1c",
          6509 => x"33575574",
          6510 => x"802ebb38",
          6511 => x"74842e09",
          6512 => x"810680e7",
          6513 => x"3875852a",
          6514 => x"70810677",
          6515 => x"822a5851",
          6516 => x"5473802e",
          6517 => x"96387581",
          6518 => x"06547380",
          6519 => x"2efbb538",
          6520 => x"ff800bab",
          6521 => x"1c348055",
          6522 => x"80c13975",
          6523 => x"81065473",
          6524 => x"ba388555",
          6525 => x"b6397582",
          6526 => x"2a708106",
          6527 => x"515473ab",
          6528 => x"38861b33",
          6529 => x"70842a70",
          6530 => x"81065155",
          6531 => x"5573802e",
          6532 => x"e138901b",
          6533 => x"0883ff06",
          6534 => x"1db40552",
          6535 => x"7c51f5db",
          6536 => x"3f82b698",
          6537 => x"08881c0c",
          6538 => x"faea3974",
          6539 => x"82b6980c",
          6540 => x"8f3d0d04",
          6541 => x"f63d0d7c",
          6542 => x"5bff7b08",
          6543 => x"70717355",
          6544 => x"595c5559",
          6545 => x"73802e81",
          6546 => x"c6387570",
          6547 => x"81055733",
          6548 => x"70a02652",
          6549 => x"5271ba2e",
          6550 => x"8d3870ee",
          6551 => x"3871ba2e",
          6552 => x"09810681",
          6553 => x"a5387333",
          6554 => x"d0117081",
          6555 => x"ff065152",
          6556 => x"53708926",
          6557 => x"91388214",
          6558 => x"7381ff06",
          6559 => x"d0055652",
          6560 => x"71762e80",
          6561 => x"f738800b",
          6562 => x"82afd059",
          6563 => x"5577087a",
          6564 => x"55577670",
          6565 => x"81055833",
          6566 => x"74708105",
          6567 => x"5633ff9f",
          6568 => x"12535353",
          6569 => x"70992689",
          6570 => x"38e01370",
          6571 => x"81ff0654",
          6572 => x"51ff9f12",
          6573 => x"51709926",
          6574 => x"8938e012",
          6575 => x"7081ff06",
          6576 => x"53517230",
          6577 => x"709f2a51",
          6578 => x"5172722e",
          6579 => x"09810685",
          6580 => x"3870ffbe",
          6581 => x"38723074",
          6582 => x"77327030",
          6583 => x"7072079f",
          6584 => x"2a739f2a",
          6585 => x"07535454",
          6586 => x"5170802e",
          6587 => x"8f388115",
          6588 => x"84195955",
          6589 => x"837525ff",
          6590 => x"94388b39",
          6591 => x"74832486",
          6592 => x"3874767c",
          6593 => x"0c597851",
          6594 => x"863982cd",
          6595 => x"e4335170",
          6596 => x"82b6980c",
          6597 => x"8c3d0d04",
          6598 => x"fa3d0d78",
          6599 => x"56800b83",
          6600 => x"1734ff0b",
          6601 => x"b0170c79",
          6602 => x"527551e2",
          6603 => x"e03f8455",
          6604 => x"82b69808",
          6605 => x"81803884",
          6606 => x"b21651df",
          6607 => x"b43f82b6",
          6608 => x"980883ff",
          6609 => x"ff065483",
          6610 => x"557382d4",
          6611 => x"d52e0981",
          6612 => x"0680e338",
          6613 => x"800bb417",
          6614 => x"33565774",
          6615 => x"81e92e09",
          6616 => x"81068338",
          6617 => x"81577481",
          6618 => x"eb327030",
          6619 => x"70802579",
          6620 => x"07515154",
          6621 => x"738a3874",
          6622 => x"81e82e09",
          6623 => x"8106b538",
          6624 => x"835382af",
          6625 => x"905280ea",
          6626 => x"1651e0b1",
          6627 => x"3f82b698",
          6628 => x"085582b6",
          6629 => x"9808802e",
          6630 => x"9d388553",
          6631 => x"82af9452",
          6632 => x"81861651",
          6633 => x"e0973f82",
          6634 => x"b6980855",
          6635 => x"82b69808",
          6636 => x"802e8338",
          6637 => x"82557482",
          6638 => x"b6980c88",
          6639 => x"3d0d04f2",
          6640 => x"3d0d6102",
          6641 => x"840580cb",
          6642 => x"05335855",
          6643 => x"80750c60",
          6644 => x"51fce13f",
          6645 => x"82b69808",
          6646 => x"588b5680",
          6647 => x"0b82b698",
          6648 => x"082486fc",
          6649 => x"3882b698",
          6650 => x"08842982",
          6651 => x"cdd00570",
          6652 => x"0855538c",
          6653 => x"5673802e",
          6654 => x"86e63873",
          6655 => x"750c7681",
          6656 => x"fe067433",
          6657 => x"54577280",
          6658 => x"2eae3881",
          6659 => x"143351d7",
          6660 => x"ca3f82b6",
          6661 => x"980881ff",
          6662 => x"06708106",
          6663 => x"54557298",
          6664 => x"3876802e",
          6665 => x"86b83874",
          6666 => x"822a7081",
          6667 => x"0651538a",
          6668 => x"567286ac",
          6669 => x"3886a739",
          6670 => x"80743477",
          6671 => x"81153481",
          6672 => x"52811433",
          6673 => x"51d7b23f",
          6674 => x"82b69808",
          6675 => x"81ff0670",
          6676 => x"81065455",
          6677 => x"83567286",
          6678 => x"87387680",
          6679 => x"2e8f3874",
          6680 => x"822a7081",
          6681 => x"0651538a",
          6682 => x"567285f4",
          6683 => x"38807053",
          6684 => x"74525bfd",
          6685 => x"a33f82b6",
          6686 => x"980881ff",
          6687 => x"06577682",
          6688 => x"2e098106",
          6689 => x"80e2388c",
          6690 => x"3d745658",
          6691 => x"835683f6",
          6692 => x"15337058",
          6693 => x"5372802e",
          6694 => x"8d3883fa",
          6695 => x"1551dce8",
          6696 => x"3f82b698",
          6697 => x"08577678",
          6698 => x"7084055a",
          6699 => x"0cff1690",
          6700 => x"16565675",
          6701 => x"8025d738",
          6702 => x"800b8d3d",
          6703 => x"54567270",
          6704 => x"84055408",
          6705 => x"5b83577a",
          6706 => x"802e9538",
          6707 => x"7a527351",
          6708 => x"fcc63f82",
          6709 => x"b6980881",
          6710 => x"ff065781",
          6711 => x"77278938",
          6712 => x"81165683",
          6713 => x"7627d738",
          6714 => x"81567684",
          6715 => x"2e84f138",
          6716 => x"8d567681",
          6717 => x"2684e938",
          6718 => x"bf1451db",
          6719 => x"f43f82b6",
          6720 => x"980883ff",
          6721 => x"ff065372",
          6722 => x"84802e09",
          6723 => x"810684d0",
          6724 => x"3880ca14",
          6725 => x"51dbda3f",
          6726 => x"82b69808",
          6727 => x"83ffff06",
          6728 => x"58778d38",
          6729 => x"80d81451",
          6730 => x"dbde3f82",
          6731 => x"b6980858",
          6732 => x"779c150c",
          6733 => x"80c41433",
          6734 => x"82153480",
          6735 => x"c41433ff",
          6736 => x"117081ff",
          6737 => x"06515455",
          6738 => x"8d567281",
          6739 => x"26849138",
          6740 => x"7481ff06",
          6741 => x"78712980",
          6742 => x"c1163352",
          6743 => x"5953728a",
          6744 => x"15237280",
          6745 => x"2e8b38ff",
          6746 => x"13730653",
          6747 => x"72802e86",
          6748 => x"388d5683",
          6749 => x"eb3980c5",
          6750 => x"1451daf5",
          6751 => x"3f82b698",
          6752 => x"085382b6",
          6753 => x"98088815",
          6754 => x"23728f06",
          6755 => x"578d5676",
          6756 => x"83ce3880",
          6757 => x"c71451da",
          6758 => x"d83f82b6",
          6759 => x"980883ff",
          6760 => x"ff065574",
          6761 => x"8d3880d4",
          6762 => x"1451dadc",
          6763 => x"3f82b698",
          6764 => x"085580c2",
          6765 => x"1451dab9",
          6766 => x"3f82b698",
          6767 => x"0883ffff",
          6768 => x"06538d56",
          6769 => x"72802e83",
          6770 => x"97388814",
          6771 => x"22781471",
          6772 => x"842a055a",
          6773 => x"5a787526",
          6774 => x"8386388a",
          6775 => x"14225274",
          6776 => x"793151fe",
          6777 => x"f39d3f82",
          6778 => x"b6980855",
          6779 => x"82b69808",
          6780 => x"802e82ec",
          6781 => x"3882b698",
          6782 => x"0880ffff",
          6783 => x"fff52683",
          6784 => x"38835774",
          6785 => x"83fff526",
          6786 => x"83388257",
          6787 => x"749ff526",
          6788 => x"85388157",
          6789 => x"89398d56",
          6790 => x"76802e82",
          6791 => x"c3388215",
          6792 => x"7098160c",
          6793 => x"7ba0160c",
          6794 => x"731c70a4",
          6795 => x"170c7a1d",
          6796 => x"ac170c54",
          6797 => x"5576832e",
          6798 => x"098106af",
          6799 => x"3880de14",
          6800 => x"51d9ae3f",
          6801 => x"82b69808",
          6802 => x"83ffff06",
          6803 => x"538d5672",
          6804 => x"828e3879",
          6805 => x"828a3880",
          6806 => x"e01451d9",
          6807 => x"ab3f82b6",
          6808 => x"9808a815",
          6809 => x"0c74822b",
          6810 => x"53a2398d",
          6811 => x"5679802e",
          6812 => x"81ee3877",
          6813 => x"13a8150c",
          6814 => x"74155376",
          6815 => x"822e8d38",
          6816 => x"74101570",
          6817 => x"812a7681",
          6818 => x"06055153",
          6819 => x"83ff1389",
          6820 => x"2a538d56",
          6821 => x"729c1508",
          6822 => x"2681c538",
          6823 => x"ff0b9015",
          6824 => x"0cff0b8c",
          6825 => x"150cff80",
          6826 => x"0b841534",
          6827 => x"76832e09",
          6828 => x"81068192",
          6829 => x"3880e414",
          6830 => x"51d8b63f",
          6831 => x"82b69808",
          6832 => x"83ffff06",
          6833 => x"5372812e",
          6834 => x"09810680",
          6835 => x"f938811b",
          6836 => x"527351db",
          6837 => x"b83f82b6",
          6838 => x"980880ea",
          6839 => x"3882b698",
          6840 => x"08841534",
          6841 => x"84b21451",
          6842 => x"d8873f82",
          6843 => x"b6980883",
          6844 => x"ffff0653",
          6845 => x"7282d4d5",
          6846 => x"2e098106",
          6847 => x"80c838b4",
          6848 => x"1451d884",
          6849 => x"3f82b698",
          6850 => x"08848b85",
          6851 => x"a4d22e09",
          6852 => x"8106b338",
          6853 => x"84981451",
          6854 => x"d7ee3f82",
          6855 => x"b6980886",
          6856 => x"8a85e4f2",
          6857 => x"2e098106",
          6858 => x"9d38849c",
          6859 => x"1451d7d8",
          6860 => x"3f82b698",
          6861 => x"0890150c",
          6862 => x"84a01451",
          6863 => x"d7ca3f82",
          6864 => x"b698088c",
          6865 => x"150c7674",
          6866 => x"3482cde0",
          6867 => x"22810553",
          6868 => x"7282cde0",
          6869 => x"23728615",
          6870 => x"23800b94",
          6871 => x"150c8056",
          6872 => x"7582b698",
          6873 => x"0c903d0d",
          6874 => x"04fb3d0d",
          6875 => x"77548955",
          6876 => x"73802eb9",
          6877 => x"38730853",
          6878 => x"72802eb1",
          6879 => x"38723352",
          6880 => x"71802ea9",
          6881 => x"38861322",
          6882 => x"84152257",
          6883 => x"5271762e",
          6884 => x"09810699",
          6885 => x"38811333",
          6886 => x"51d0c03f",
          6887 => x"82b69808",
          6888 => x"81065271",
          6889 => x"88387174",
          6890 => x"08545583",
          6891 => x"39805378",
          6892 => x"73710c52",
          6893 => x"7482b698",
          6894 => x"0c873d0d",
          6895 => x"04fa3d0d",
          6896 => x"02ab0533",
          6897 => x"7a58893d",
          6898 => x"fc055256",
          6899 => x"f4e63f8b",
          6900 => x"54800b82",
          6901 => x"b6980824",
          6902 => x"bc3882b6",
          6903 => x"98088429",
          6904 => x"82cdd005",
          6905 => x"70085555",
          6906 => x"73802e84",
          6907 => x"38807434",
          6908 => x"78547380",
          6909 => x"2e843880",
          6910 => x"74347875",
          6911 => x"0c755475",
          6912 => x"802e9238",
          6913 => x"8053893d",
          6914 => x"70538405",
          6915 => x"51f7b03f",
          6916 => x"82b69808",
          6917 => x"547382b6",
          6918 => x"980c883d",
          6919 => x"0d04eb3d",
          6920 => x"0d670284",
          6921 => x"0580e705",
          6922 => x"33595989",
          6923 => x"5478802e",
          6924 => x"84c83877",
          6925 => x"bf067054",
          6926 => x"983dd005",
          6927 => x"53993d84",
          6928 => x"055258f6",
          6929 => x"fa3f82b6",
          6930 => x"98085582",
          6931 => x"b6980884",
          6932 => x"a4387a5c",
          6933 => x"68528c3d",
          6934 => x"705256ed",
          6935 => x"c63f82b6",
          6936 => x"98085582",
          6937 => x"b6980892",
          6938 => x"380280d7",
          6939 => x"05337098",
          6940 => x"2b555773",
          6941 => x"80258338",
          6942 => x"8655779c",
          6943 => x"06547380",
          6944 => x"2e81ab38",
          6945 => x"74802e95",
          6946 => x"3874842e",
          6947 => x"098106aa",
          6948 => x"387551ea",
          6949 => x"f83f82b6",
          6950 => x"9808559e",
          6951 => x"3902b205",
          6952 => x"33910654",
          6953 => x"7381b838",
          6954 => x"77822a70",
          6955 => x"81065154",
          6956 => x"73802e8e",
          6957 => x"38885583",
          6958 => x"bc397788",
          6959 => x"07587483",
          6960 => x"b4387783",
          6961 => x"2a708106",
          6962 => x"51547380",
          6963 => x"2e81af38",
          6964 => x"62527a51",
          6965 => x"e8a53f82",
          6966 => x"b6980856",
          6967 => x"8288b20a",
          6968 => x"52628e05",
          6969 => x"51d4ea3f",
          6970 => x"6254a00b",
          6971 => x"8b153480",
          6972 => x"5362527a",
          6973 => x"51e8bd3f",
          6974 => x"8052629c",
          6975 => x"0551d4d1",
          6976 => x"3f7a5481",
          6977 => x"0b831534",
          6978 => x"75802e80",
          6979 => x"f1387ab0",
          6980 => x"11085154",
          6981 => x"80537552",
          6982 => x"973dd405",
          6983 => x"51ddbe3f",
          6984 => x"82b69808",
          6985 => x"5582b698",
          6986 => x"0882ca38",
          6987 => x"b7397482",
          6988 => x"c43802b2",
          6989 => x"05337084",
          6990 => x"2a708106",
          6991 => x"51555673",
          6992 => x"802e8638",
          6993 => x"845582ad",
          6994 => x"3977812a",
          6995 => x"70810651",
          6996 => x"5473802e",
          6997 => x"a9387581",
          6998 => x"06547380",
          6999 => x"2ea03887",
          7000 => x"55829239",
          7001 => x"73527a51",
          7002 => x"d6a33f82",
          7003 => x"b698087b",
          7004 => x"ff188c12",
          7005 => x"0c555582",
          7006 => x"b6980881",
          7007 => x"f8387783",
          7008 => x"2a708106",
          7009 => x"51547380",
          7010 => x"2e863877",
          7011 => x"80c00758",
          7012 => x"7ab01108",
          7013 => x"a01b0c63",
          7014 => x"a41b0c63",
          7015 => x"53705257",
          7016 => x"e6d93f82",
          7017 => x"b6980882",
          7018 => x"b6980888",
          7019 => x"1b0c639c",
          7020 => x"05525ad2",
          7021 => x"d33f82b6",
          7022 => x"980882b6",
          7023 => x"98088c1b",
          7024 => x"0c777a0c",
          7025 => x"56861722",
          7026 => x"841a2377",
          7027 => x"901a3480",
          7028 => x"0b911a34",
          7029 => x"800b9c1a",
          7030 => x"0c800b94",
          7031 => x"1a0c7785",
          7032 => x"2a708106",
          7033 => x"51547380",
          7034 => x"2e818d38",
          7035 => x"82b69808",
          7036 => x"802e8184",
          7037 => x"3882b698",
          7038 => x"08941a0c",
          7039 => x"8a172270",
          7040 => x"892b7b52",
          7041 => x"5957a839",
          7042 => x"76527851",
          7043 => x"d79f3f82",
          7044 => x"b6980857",
          7045 => x"82b69808",
          7046 => x"81268338",
          7047 => x"825582b6",
          7048 => x"9808ff2e",
          7049 => x"09810683",
          7050 => x"38795575",
          7051 => x"78315674",
          7052 => x"30707607",
          7053 => x"80255154",
          7054 => x"7776278a",
          7055 => x"38817075",
          7056 => x"06555a73",
          7057 => x"c3387698",
          7058 => x"1a0c74a9",
          7059 => x"387583ff",
          7060 => x"06547380",
          7061 => x"2ea23876",
          7062 => x"527a51d6",
          7063 => x"a63f82b6",
          7064 => x"98088538",
          7065 => x"82558e39",
          7066 => x"75892a82",
          7067 => x"b6980805",
          7068 => x"9c1a0c84",
          7069 => x"3980790c",
          7070 => x"74547382",
          7071 => x"b6980c97",
          7072 => x"3d0d04f2",
          7073 => x"3d0d6063",
          7074 => x"65644040",
          7075 => x"5d59807e",
          7076 => x"0c903dfc",
          7077 => x"05527851",
          7078 => x"f9cf3f82",
          7079 => x"b6980855",
          7080 => x"82b69808",
          7081 => x"8a389119",
          7082 => x"33557480",
          7083 => x"2e863874",
          7084 => x"5682c439",
          7085 => x"90193381",
          7086 => x"06558756",
          7087 => x"74802e82",
          7088 => x"b6389539",
          7089 => x"820b911a",
          7090 => x"34825682",
          7091 => x"aa39810b",
          7092 => x"911a3481",
          7093 => x"5682a039",
          7094 => x"8c190894",
          7095 => x"1a083155",
          7096 => x"747c2783",
          7097 => x"38745c7b",
          7098 => x"802e8289",
          7099 => x"38941908",
          7100 => x"7083ff06",
          7101 => x"56567481",
          7102 => x"b2387e8a",
          7103 => x"1122ff05",
          7104 => x"77892a06",
          7105 => x"5b5579a8",
          7106 => x"38758738",
          7107 => x"88190855",
          7108 => x"8f399819",
          7109 => x"08527851",
          7110 => x"d5933f82",
          7111 => x"b6980855",
          7112 => x"817527ff",
          7113 => x"9f3874ff",
          7114 => x"2effa338",
          7115 => x"74981a0c",
          7116 => x"98190852",
          7117 => x"7e51d4cb",
          7118 => x"3f82b698",
          7119 => x"08802eff",
          7120 => x"833882b6",
          7121 => x"98081a7c",
          7122 => x"892a5957",
          7123 => x"77802e80",
          7124 => x"d638771a",
          7125 => x"7f8a1122",
          7126 => x"585c5575",
          7127 => x"75278538",
          7128 => x"757a3158",
          7129 => x"77547653",
          7130 => x"7c52811b",
          7131 => x"3351ca88",
          7132 => x"3f82b698",
          7133 => x"08fed738",
          7134 => x"7e831133",
          7135 => x"56567480",
          7136 => x"2e9f38b0",
          7137 => x"16087731",
          7138 => x"55747827",
          7139 => x"94388480",
          7140 => x"53b41652",
          7141 => x"b0160877",
          7142 => x"31892b7d",
          7143 => x"0551cfe0",
          7144 => x"3f77892b",
          7145 => x"56b93976",
          7146 => x"9c1a0c94",
          7147 => x"190883ff",
          7148 => x"06848071",
          7149 => x"3157557b",
          7150 => x"76278338",
          7151 => x"7b569c19",
          7152 => x"08527e51",
          7153 => x"d1c73f82",
          7154 => x"b69808fe",
          7155 => x"81387553",
          7156 => x"94190883",
          7157 => x"ff061fb4",
          7158 => x"05527c51",
          7159 => x"cfa23f7b",
          7160 => x"76317e08",
          7161 => x"177f0c76",
          7162 => x"1e941b08",
          7163 => x"18941c0c",
          7164 => x"5e5cfdf3",
          7165 => x"39805675",
          7166 => x"82b6980c",
          7167 => x"903d0d04",
          7168 => x"f23d0d60",
          7169 => x"63656440",
          7170 => x"405d5880",
          7171 => x"7e0c903d",
          7172 => x"fc055277",
          7173 => x"51f6d23f",
          7174 => x"82b69808",
          7175 => x"5582b698",
          7176 => x"088a3891",
          7177 => x"18335574",
          7178 => x"802e8638",
          7179 => x"745683b8",
          7180 => x"39901833",
          7181 => x"70812a70",
          7182 => x"81065156",
          7183 => x"56875674",
          7184 => x"802e83a4",
          7185 => x"38953982",
          7186 => x"0b911934",
          7187 => x"82568398",
          7188 => x"39810b91",
          7189 => x"19348156",
          7190 => x"838e3994",
          7191 => x"18087c11",
          7192 => x"56567476",
          7193 => x"27843875",
          7194 => x"095c7b80",
          7195 => x"2e82ec38",
          7196 => x"94180870",
          7197 => x"83ff0656",
          7198 => x"567481fd",
          7199 => x"387e8a11",
          7200 => x"22ff0577",
          7201 => x"892a065c",
          7202 => x"557abf38",
          7203 => x"758c3888",
          7204 => x"18085574",
          7205 => x"9c387a52",
          7206 => x"85399818",
          7207 => x"08527751",
          7208 => x"d7e73f82",
          7209 => x"b6980855",
          7210 => x"82b69808",
          7211 => x"802e82ab",
          7212 => x"3874812e",
          7213 => x"ff913874",
          7214 => x"ff2eff95",
          7215 => x"38749819",
          7216 => x"0c881808",
          7217 => x"85387488",
          7218 => x"190c7e55",
          7219 => x"b015089c",
          7220 => x"19082e09",
          7221 => x"81068d38",
          7222 => x"7451cec1",
          7223 => x"3f82b698",
          7224 => x"08feee38",
          7225 => x"98180852",
          7226 => x"7e51d197",
          7227 => x"3f82b698",
          7228 => x"08802efe",
          7229 => x"d23882b6",
          7230 => x"98081b7c",
          7231 => x"892a5a57",
          7232 => x"78802e80",
          7233 => x"d538781b",
          7234 => x"7f8a1122",
          7235 => x"585b5575",
          7236 => x"75278538",
          7237 => x"757b3159",
          7238 => x"78547653",
          7239 => x"7c52811a",
          7240 => x"3351c8be",
          7241 => x"3f82b698",
          7242 => x"08fea638",
          7243 => x"7eb01108",
          7244 => x"78315656",
          7245 => x"7479279b",
          7246 => x"38848053",
          7247 => x"b0160877",
          7248 => x"31892b7d",
          7249 => x"0552b416",
          7250 => x"51ccb53f",
          7251 => x"7e55800b",
          7252 => x"83163478",
          7253 => x"892b5680",
          7254 => x"db398c18",
          7255 => x"08941908",
          7256 => x"2693387e",
          7257 => x"51cdb63f",
          7258 => x"82b69808",
          7259 => x"fde3387e",
          7260 => x"77b0120c",
          7261 => x"55769c19",
          7262 => x"0c941808",
          7263 => x"83ff0684",
          7264 => x"80713157",
          7265 => x"557b7627",
          7266 => x"83387b56",
          7267 => x"9c180852",
          7268 => x"7e51cdf9",
          7269 => x"3f82b698",
          7270 => x"08fdb638",
          7271 => x"75537c52",
          7272 => x"94180883",
          7273 => x"ff061fb4",
          7274 => x"0551cbd4",
          7275 => x"3f7e5581",
          7276 => x"0b831634",
          7277 => x"7b76317e",
          7278 => x"08177f0c",
          7279 => x"761e941a",
          7280 => x"08187094",
          7281 => x"1c0c8c1b",
          7282 => x"0858585e",
          7283 => x"5c747627",
          7284 => x"83387555",
          7285 => x"748c190c",
          7286 => x"fd903990",
          7287 => x"183380c0",
          7288 => x"07557490",
          7289 => x"19348056",
          7290 => x"7582b698",
          7291 => x"0c903d0d",
          7292 => x"04f83d0d",
          7293 => x"7a8b3dfc",
          7294 => x"05537052",
          7295 => x"56f2ea3f",
          7296 => x"82b69808",
          7297 => x"5782b698",
          7298 => x"0880fb38",
          7299 => x"90163370",
          7300 => x"862a7081",
          7301 => x"06515555",
          7302 => x"73802e80",
          7303 => x"e938a016",
          7304 => x"08527851",
          7305 => x"cce73f82",
          7306 => x"b6980857",
          7307 => x"82b69808",
          7308 => x"80d438a4",
          7309 => x"16088b11",
          7310 => x"33a00755",
          7311 => x"55738b16",
          7312 => x"34881608",
          7313 => x"53745275",
          7314 => x"0851dde8",
          7315 => x"3f8c1608",
          7316 => x"529c1551",
          7317 => x"c9fb3f82",
          7318 => x"88b20a52",
          7319 => x"961551c9",
          7320 => x"f03f7652",
          7321 => x"921551c9",
          7322 => x"ca3f7854",
          7323 => x"810b8315",
          7324 => x"347851cc",
          7325 => x"df3f82b6",
          7326 => x"98089017",
          7327 => x"3381bf06",
          7328 => x"55577390",
          7329 => x"17347682",
          7330 => x"b6980c8a",
          7331 => x"3d0d04fc",
          7332 => x"3d0d7670",
          7333 => x"5254fed9",
          7334 => x"3f82b698",
          7335 => x"085382b6",
          7336 => x"98089c38",
          7337 => x"863dfc05",
          7338 => x"527351f1",
          7339 => x"bc3f82b6",
          7340 => x"98085382",
          7341 => x"b6980887",
          7342 => x"3882b698",
          7343 => x"08740c72",
          7344 => x"82b6980c",
          7345 => x"863d0d04",
          7346 => x"ff3d0d84",
          7347 => x"3d51e6e4",
          7348 => x"3f8b5280",
          7349 => x"0b82b698",
          7350 => x"08248b38",
          7351 => x"82b69808",
          7352 => x"82cde434",
          7353 => x"80527182",
          7354 => x"b6980c83",
          7355 => x"3d0d04ef",
          7356 => x"3d0d8053",
          7357 => x"933dd005",
          7358 => x"52943d51",
          7359 => x"e9c13f82",
          7360 => x"b6980855",
          7361 => x"82b69808",
          7362 => x"80e03876",
          7363 => x"58635293",
          7364 => x"3dd40551",
          7365 => x"e08d3f82",
          7366 => x"b6980855",
          7367 => x"82b69808",
          7368 => x"bc380280",
          7369 => x"c7053370",
          7370 => x"982b5556",
          7371 => x"73802589",
          7372 => x"38767a94",
          7373 => x"120c54b2",
          7374 => x"3902a205",
          7375 => x"3370842a",
          7376 => x"70810651",
          7377 => x"55567380",
          7378 => x"2e9e3876",
          7379 => x"7f537052",
          7380 => x"54dba83f",
          7381 => x"82b69808",
          7382 => x"94150c8e",
          7383 => x"3982b698",
          7384 => x"08842e09",
          7385 => x"81068338",
          7386 => x"85557482",
          7387 => x"b6980c93",
          7388 => x"3d0d04e4",
          7389 => x"3d0d6f6f",
          7390 => x"5b5b807a",
          7391 => x"3480539e",
          7392 => x"3dffb805",
          7393 => x"529f3d51",
          7394 => x"e8b53f82",
          7395 => x"b6980857",
          7396 => x"82b69808",
          7397 => x"82fc387b",
          7398 => x"437a7c94",
          7399 => x"11084755",
          7400 => x"58645473",
          7401 => x"802e81ed",
          7402 => x"38a05293",
          7403 => x"3d705255",
          7404 => x"d5ea3f82",
          7405 => x"b6980857",
          7406 => x"82b69808",
          7407 => x"82d43868",
          7408 => x"527b51c9",
          7409 => x"c83f82b6",
          7410 => x"98085782",
          7411 => x"b6980882",
          7412 => x"c1386952",
          7413 => x"7b51daa3",
          7414 => x"3f82b698",
          7415 => x"08457652",
          7416 => x"7451d5b8",
          7417 => x"3f82b698",
          7418 => x"085782b6",
          7419 => x"980882a2",
          7420 => x"38805274",
          7421 => x"51daeb3f",
          7422 => x"82b69808",
          7423 => x"5782b698",
          7424 => x"08a43869",
          7425 => x"527b51d9",
          7426 => x"f23f7382",
          7427 => x"b698082e",
          7428 => x"a6387652",
          7429 => x"7451d6cf",
          7430 => x"3f82b698",
          7431 => x"085782b6",
          7432 => x"9808802e",
          7433 => x"cc387684",
          7434 => x"2e098106",
          7435 => x"86388257",
          7436 => x"81e03976",
          7437 => x"81dc389e",
          7438 => x"3dffbc05",
          7439 => x"527451dc",
          7440 => x"c93f7690",
          7441 => x"3d781181",
          7442 => x"11335156",
          7443 => x"5a567380",
          7444 => x"2e913802",
          7445 => x"b9055581",
          7446 => x"16811670",
          7447 => x"33565656",
          7448 => x"73f53881",
          7449 => x"16547378",
          7450 => x"26819038",
          7451 => x"75802e99",
          7452 => x"38781681",
          7453 => x"0555ff18",
          7454 => x"6f11ff18",
          7455 => x"ff185858",
          7456 => x"55587433",
          7457 => x"743475ee",
          7458 => x"38ff186f",
          7459 => x"115558af",
          7460 => x"7434fe8d",
          7461 => x"39777b2e",
          7462 => x"0981068a",
          7463 => x"38ff186f",
          7464 => x"115558af",
          7465 => x"7434800b",
          7466 => x"82cde433",
          7467 => x"70842982",
          7468 => x"afd00570",
          7469 => x"08703352",
          7470 => x"5c565656",
          7471 => x"73762e8d",
          7472 => x"38811670",
          7473 => x"1a703351",
          7474 => x"555673f5",
          7475 => x"38821654",
          7476 => x"737826a7",
          7477 => x"38805574",
          7478 => x"76279138",
          7479 => x"74195473",
          7480 => x"337a7081",
          7481 => x"055c3481",
          7482 => x"1555ec39",
          7483 => x"ba7a7081",
          7484 => x"055c3474",
          7485 => x"ff2e0981",
          7486 => x"06853891",
          7487 => x"5794396e",
          7488 => x"18811959",
          7489 => x"5473337a",
          7490 => x"7081055c",
          7491 => x"347a7826",
          7492 => x"ee38807a",
          7493 => x"347682b6",
          7494 => x"980c9e3d",
          7495 => x"0d04f73d",
          7496 => x"0d7b7d8d",
          7497 => x"3dfc0554",
          7498 => x"71535755",
          7499 => x"ecbb3f82",
          7500 => x"b6980853",
          7501 => x"82b69808",
          7502 => x"82fa3891",
          7503 => x"15335372",
          7504 => x"82f2388c",
          7505 => x"15085473",
          7506 => x"76279238",
          7507 => x"90153370",
          7508 => x"812a7081",
          7509 => x"06515457",
          7510 => x"72833873",
          7511 => x"56941508",
          7512 => x"54807094",
          7513 => x"170c5875",
          7514 => x"782e8297",
          7515 => x"38798a11",
          7516 => x"2270892b",
          7517 => x"59515373",
          7518 => x"782eb738",
          7519 => x"7652ff16",
          7520 => x"51fedbff",
          7521 => x"3f82b698",
          7522 => x"08ff1578",
          7523 => x"54705355",
          7524 => x"53fedbef",
          7525 => x"3f82b698",
          7526 => x"08732696",
          7527 => x"38763070",
          7528 => x"75067094",
          7529 => x"180c7771",
          7530 => x"31981808",
          7531 => x"57585153",
          7532 => x"b1398815",
          7533 => x"085473a6",
          7534 => x"38735274",
          7535 => x"51cdca3f",
          7536 => x"82b69808",
          7537 => x"5482b698",
          7538 => x"08812e81",
          7539 => x"9a3882b6",
          7540 => x"9808ff2e",
          7541 => x"819b3882",
          7542 => x"b6980888",
          7543 => x"160c7398",
          7544 => x"160c7380",
          7545 => x"2e819c38",
          7546 => x"76762780",
          7547 => x"dc387577",
          7548 => x"31941608",
          7549 => x"1894170c",
          7550 => x"90163370",
          7551 => x"812a7081",
          7552 => x"0651555a",
          7553 => x"5672802e",
          7554 => x"9a387352",
          7555 => x"7451ccf9",
          7556 => x"3f82b698",
          7557 => x"085482b6",
          7558 => x"98089438",
          7559 => x"82b69808",
          7560 => x"56a73973",
          7561 => x"527451c7",
          7562 => x"843f82b6",
          7563 => x"98085473",
          7564 => x"ff2ebe38",
          7565 => x"817427af",
          7566 => x"38795373",
          7567 => x"98140827",
          7568 => x"a6387398",
          7569 => x"160cffa0",
          7570 => x"39941508",
          7571 => x"1694160c",
          7572 => x"7583ff06",
          7573 => x"5372802e",
          7574 => x"aa387352",
          7575 => x"7951c6a3",
          7576 => x"3f82b698",
          7577 => x"08943882",
          7578 => x"0b911634",
          7579 => x"825380c4",
          7580 => x"39810b91",
          7581 => x"16348153",
          7582 => x"bb397589",
          7583 => x"2a82b698",
          7584 => x"08055894",
          7585 => x"1508548c",
          7586 => x"15087427",
          7587 => x"9038738c",
          7588 => x"160c9015",
          7589 => x"3380c007",
          7590 => x"53729016",
          7591 => x"347383ff",
          7592 => x"06537280",
          7593 => x"2e8c3877",
          7594 => x"9c16082e",
          7595 => x"8538779c",
          7596 => x"160c8053",
          7597 => x"7282b698",
          7598 => x"0c8b3d0d",
          7599 => x"04f93d0d",
          7600 => x"79568954",
          7601 => x"75802e81",
          7602 => x"8a388053",
          7603 => x"893dfc05",
          7604 => x"528a3d84",
          7605 => x"0551e1e7",
          7606 => x"3f82b698",
          7607 => x"085582b6",
          7608 => x"980880ea",
          7609 => x"3877760c",
          7610 => x"7a527551",
          7611 => x"d8b53f82",
          7612 => x"b6980855",
          7613 => x"82b69808",
          7614 => x"80c338ab",
          7615 => x"16337098",
          7616 => x"2b555780",
          7617 => x"7424a238",
          7618 => x"86163370",
          7619 => x"842a7081",
          7620 => x"06515557",
          7621 => x"73802ead",
          7622 => x"389c1608",
          7623 => x"527751d3",
          7624 => x"da3f82b6",
          7625 => x"98088817",
          7626 => x"0c775486",
          7627 => x"14228417",
          7628 => x"23745275",
          7629 => x"51cee53f",
          7630 => x"82b69808",
          7631 => x"5574842e",
          7632 => x"09810685",
          7633 => x"38855586",
          7634 => x"3974802e",
          7635 => x"84388076",
          7636 => x"0c745473",
          7637 => x"82b6980c",
          7638 => x"893d0d04",
          7639 => x"fc3d0d76",
          7640 => x"873dfc05",
          7641 => x"53705253",
          7642 => x"e7ff3f82",
          7643 => x"b6980887",
          7644 => x"3882b698",
          7645 => x"08730c86",
          7646 => x"3d0d04fb",
          7647 => x"3d0d7779",
          7648 => x"893dfc05",
          7649 => x"54715356",
          7650 => x"54e7de3f",
          7651 => x"82b69808",
          7652 => x"5382b698",
          7653 => x"0880df38",
          7654 => x"74933882",
          7655 => x"b6980852",
          7656 => x"7351cdf8",
          7657 => x"3f82b698",
          7658 => x"085380ca",
          7659 => x"3982b698",
          7660 => x"08527351",
          7661 => x"d3ac3f82",
          7662 => x"b6980853",
          7663 => x"82b69808",
          7664 => x"842e0981",
          7665 => x"06853880",
          7666 => x"53873982",
          7667 => x"b69808a6",
          7668 => x"38745273",
          7669 => x"51d5b33f",
          7670 => x"72527351",
          7671 => x"cf893f82",
          7672 => x"b6980884",
          7673 => x"32703070",
          7674 => x"72079f2c",
          7675 => x"7082b698",
          7676 => x"08065151",
          7677 => x"54547282",
          7678 => x"b6980c87",
          7679 => x"3d0d04ee",
          7680 => x"3d0d6557",
          7681 => x"8053893d",
          7682 => x"7053963d",
          7683 => x"5256dfaf",
          7684 => x"3f82b698",
          7685 => x"085582b6",
          7686 => x"9808b238",
          7687 => x"64527551",
          7688 => x"d6813f82",
          7689 => x"b6980855",
          7690 => x"82b69808",
          7691 => x"a0380280",
          7692 => x"cb053370",
          7693 => x"982b5558",
          7694 => x"73802585",
          7695 => x"3886558d",
          7696 => x"3976802e",
          7697 => x"88387652",
          7698 => x"7551d4be",
          7699 => x"3f7482b6",
          7700 => x"980c943d",
          7701 => x"0d04f03d",
          7702 => x"0d636555",
          7703 => x"5c805392",
          7704 => x"3dec0552",
          7705 => x"933d51de",
          7706 => x"d63f82b6",
          7707 => x"98085b82",
          7708 => x"b6980882",
          7709 => x"80387c74",
          7710 => x"0c730898",
          7711 => x"1108fe11",
          7712 => x"90130859",
          7713 => x"56585575",
          7714 => x"74269138",
          7715 => x"757c0c81",
          7716 => x"e439815b",
          7717 => x"81cc3982",
          7718 => x"5b81c739",
          7719 => x"82b69808",
          7720 => x"75335559",
          7721 => x"73812e09",
          7722 => x"8106bf38",
          7723 => x"82755f57",
          7724 => x"7652923d",
          7725 => x"f00551c1",
          7726 => x"f43f82b6",
          7727 => x"9808ff2e",
          7728 => x"d13882b6",
          7729 => x"9808812e",
          7730 => x"ce3882b6",
          7731 => x"98083070",
          7732 => x"82b69808",
          7733 => x"0780257a",
          7734 => x"0581197f",
          7735 => x"53595a54",
          7736 => x"98140877",
          7737 => x"26ca3880",
          7738 => x"f939a415",
          7739 => x"0882b698",
          7740 => x"08575875",
          7741 => x"98387752",
          7742 => x"81187d52",
          7743 => x"58ffbf8d",
          7744 => x"3f82b698",
          7745 => x"085b82b6",
          7746 => x"980880d6",
          7747 => x"387c7033",
          7748 => x"7712ff1a",
          7749 => x"5d525654",
          7750 => x"74822e09",
          7751 => x"81069e38",
          7752 => x"b41451ff",
          7753 => x"bbcb3f82",
          7754 => x"b6980883",
          7755 => x"ffff0670",
          7756 => x"30708025",
          7757 => x"1b821959",
          7758 => x"5b51549b",
          7759 => x"39b41451",
          7760 => x"ffbbc53f",
          7761 => x"82b69808",
          7762 => x"f00a0670",
          7763 => x"30708025",
          7764 => x"1b841959",
          7765 => x"5b515475",
          7766 => x"83ff067a",
          7767 => x"585679ff",
          7768 => x"9238787c",
          7769 => x"0c7c7990",
          7770 => x"120c8411",
          7771 => x"33810756",
          7772 => x"54748415",
          7773 => x"347a82b6",
          7774 => x"980c923d",
          7775 => x"0d04f93d",
          7776 => x"0d798a3d",
          7777 => x"fc055370",
          7778 => x"5257e3dd",
          7779 => x"3f82b698",
          7780 => x"085682b6",
          7781 => x"980881a8",
          7782 => x"38911733",
          7783 => x"567581a0",
          7784 => x"38901733",
          7785 => x"70812a70",
          7786 => x"81065155",
          7787 => x"55875573",
          7788 => x"802e818e",
          7789 => x"38941708",
          7790 => x"54738c18",
          7791 => x"08278180",
          7792 => x"38739b38",
          7793 => x"82b69808",
          7794 => x"53881708",
          7795 => x"527651c4",
          7796 => x"8c3f82b6",
          7797 => x"98087488",
          7798 => x"190c5680",
          7799 => x"c9399817",
          7800 => x"08527651",
          7801 => x"ffbfc63f",
          7802 => x"82b69808",
          7803 => x"ff2e0981",
          7804 => x"06833881",
          7805 => x"5682b698",
          7806 => x"08812e09",
          7807 => x"81068538",
          7808 => x"8256a339",
          7809 => x"75a03877",
          7810 => x"5482b698",
          7811 => x"08981508",
          7812 => x"27943898",
          7813 => x"17085382",
          7814 => x"b6980852",
          7815 => x"7651c3bd",
          7816 => x"3f82b698",
          7817 => x"08569417",
          7818 => x"088c180c",
          7819 => x"90173380",
          7820 => x"c0075473",
          7821 => x"90183475",
          7822 => x"802e8538",
          7823 => x"75911834",
          7824 => x"75557482",
          7825 => x"b6980c89",
          7826 => x"3d0d04e2",
          7827 => x"3d0d8253",
          7828 => x"a03dffa4",
          7829 => x"0552a13d",
          7830 => x"51dae43f",
          7831 => x"82b69808",
          7832 => x"5582b698",
          7833 => x"0881f538",
          7834 => x"7845a13d",
          7835 => x"0852953d",
          7836 => x"705258d1",
          7837 => x"ae3f82b6",
          7838 => x"98085582",
          7839 => x"b6980881",
          7840 => x"db380280",
          7841 => x"fb053370",
          7842 => x"852a7081",
          7843 => x"06515556",
          7844 => x"86557381",
          7845 => x"c7387598",
          7846 => x"2b548074",
          7847 => x"2481bd38",
          7848 => x"0280d605",
          7849 => x"33708106",
          7850 => x"58548755",
          7851 => x"7681ad38",
          7852 => x"6b527851",
          7853 => x"ccc53f82",
          7854 => x"b6980874",
          7855 => x"842a7081",
          7856 => x"06515556",
          7857 => x"73802e80",
          7858 => x"d4387854",
          7859 => x"82b69808",
          7860 => x"9415082e",
          7861 => x"81863873",
          7862 => x"5a82b698",
          7863 => x"085c7652",
          7864 => x"8a3d7052",
          7865 => x"54c7b53f",
          7866 => x"82b69808",
          7867 => x"5582b698",
          7868 => x"0880e938",
          7869 => x"82b69808",
          7870 => x"527351cc",
          7871 => x"e53f82b6",
          7872 => x"98085582",
          7873 => x"b6980886",
          7874 => x"38875580",
          7875 => x"cf3982b6",
          7876 => x"9808842e",
          7877 => x"883882b6",
          7878 => x"980880c0",
          7879 => x"387751ce",
          7880 => x"c23f82b6",
          7881 => x"980882b6",
          7882 => x"98083070",
          7883 => x"82b69808",
          7884 => x"07802551",
          7885 => x"55557580",
          7886 => x"2e943873",
          7887 => x"802e8f38",
          7888 => x"80537552",
          7889 => x"7751c195",
          7890 => x"3f82b698",
          7891 => x"0855748c",
          7892 => x"387851ff",
          7893 => x"bafe3f82",
          7894 => x"b6980855",
          7895 => x"7482b698",
          7896 => x"0ca03d0d",
          7897 => x"04e93d0d",
          7898 => x"8253993d",
          7899 => x"c005529a",
          7900 => x"3d51d8cb",
          7901 => x"3f82b698",
          7902 => x"085482b6",
          7903 => x"980882b0",
          7904 => x"38785e69",
          7905 => x"528e3d70",
          7906 => x"5258cf97",
          7907 => x"3f82b698",
          7908 => x"085482b6",
          7909 => x"98088638",
          7910 => x"88548294",
          7911 => x"3982b698",
          7912 => x"08842e09",
          7913 => x"81068288",
          7914 => x"380280df",
          7915 => x"05337085",
          7916 => x"2a810651",
          7917 => x"55865474",
          7918 => x"81f63878",
          7919 => x"5a74528a",
          7920 => x"3d705257",
          7921 => x"c1c33f82",
          7922 => x"b6980875",
          7923 => x"555682b6",
          7924 => x"98088338",
          7925 => x"875482b6",
          7926 => x"9808812e",
          7927 => x"09810683",
          7928 => x"38825482",
          7929 => x"b69808ff",
          7930 => x"2e098106",
          7931 => x"86388154",
          7932 => x"81b43973",
          7933 => x"81b03882",
          7934 => x"b6980852",
          7935 => x"7851c4a4",
          7936 => x"3f82b698",
          7937 => x"085482b6",
          7938 => x"9808819a",
          7939 => x"388b53a0",
          7940 => x"52b41951",
          7941 => x"ffb78c3f",
          7942 => x"7854ae0b",
          7943 => x"b4153478",
          7944 => x"54900bbf",
          7945 => x"15348288",
          7946 => x"b20a5280",
          7947 => x"ca1951ff",
          7948 => x"b69f3f75",
          7949 => x"5378b411",
          7950 => x"5351c9f8",
          7951 => x"3fa05378",
          7952 => x"b4115380",
          7953 => x"d40551ff",
          7954 => x"b6b63f78",
          7955 => x"54ae0b80",
          7956 => x"d515347f",
          7957 => x"537880d4",
          7958 => x"115351c9",
          7959 => x"d73f7854",
          7960 => x"810b8315",
          7961 => x"347751cb",
          7962 => x"a43f82b6",
          7963 => x"98085482",
          7964 => x"b69808b2",
          7965 => x"388288b2",
          7966 => x"0a526496",
          7967 => x"0551ffb5",
          7968 => x"d03f7553",
          7969 => x"64527851",
          7970 => x"c9aa3f64",
          7971 => x"54900b8b",
          7972 => x"15347854",
          7973 => x"810b8315",
          7974 => x"347851ff",
          7975 => x"b8b63f82",
          7976 => x"b6980854",
          7977 => x"8b398053",
          7978 => x"75527651",
          7979 => x"ffbeae3f",
          7980 => x"7382b698",
          7981 => x"0c993d0d",
          7982 => x"04da3d0d",
          7983 => x"a93d8405",
          7984 => x"51d2f13f",
          7985 => x"8253a83d",
          7986 => x"ff840552",
          7987 => x"a93d51d5",
          7988 => x"ee3f82b6",
          7989 => x"98085582",
          7990 => x"b6980882",
          7991 => x"d338784d",
          7992 => x"a93d0852",
          7993 => x"9d3d7052",
          7994 => x"58ccb83f",
          7995 => x"82b69808",
          7996 => x"5582b698",
          7997 => x"0882b938",
          7998 => x"02819b05",
          7999 => x"3381a006",
          8000 => x"54865573",
          8001 => x"82aa38a0",
          8002 => x"53a43d08",
          8003 => x"52a83dff",
          8004 => x"880551ff",
          8005 => x"b4ea3fac",
          8006 => x"53775292",
          8007 => x"3d705254",
          8008 => x"ffb4dd3f",
          8009 => x"aa3d0852",
          8010 => x"7351cbf7",
          8011 => x"3f82b698",
          8012 => x"085582b6",
          8013 => x"98089538",
          8014 => x"636f2e09",
          8015 => x"81068838",
          8016 => x"65a23d08",
          8017 => x"2e923888",
          8018 => x"5581e539",
          8019 => x"82b69808",
          8020 => x"842e0981",
          8021 => x"0681b838",
          8022 => x"7351c9b1",
          8023 => x"3f82b698",
          8024 => x"085582b6",
          8025 => x"980881c8",
          8026 => x"38685693",
          8027 => x"53a83dff",
          8028 => x"9505528d",
          8029 => x"1651ffb4",
          8030 => x"873f02af",
          8031 => x"05338b17",
          8032 => x"348b1633",
          8033 => x"70842a70",
          8034 => x"81065155",
          8035 => x"55738938",
          8036 => x"74a00754",
          8037 => x"738b1734",
          8038 => x"7854810b",
          8039 => x"8315348b",
          8040 => x"16337084",
          8041 => x"2a708106",
          8042 => x"51555573",
          8043 => x"802e80e5",
          8044 => x"386e642e",
          8045 => x"80df3875",
          8046 => x"527851c6",
          8047 => x"be3f82b6",
          8048 => x"98085278",
          8049 => x"51ffb7bb",
          8050 => x"3f825582",
          8051 => x"b6980880",
          8052 => x"2e80dd38",
          8053 => x"82b69808",
          8054 => x"527851ff",
          8055 => x"b5af3f82",
          8056 => x"b6980879",
          8057 => x"80d41158",
          8058 => x"585582b6",
          8059 => x"980880c0",
          8060 => x"38811633",
          8061 => x"5473ae2e",
          8062 => x"09810699",
          8063 => x"38635375",
          8064 => x"527651c6",
          8065 => x"af3f7854",
          8066 => x"810b8315",
          8067 => x"34873982",
          8068 => x"b698089c",
          8069 => x"387751c8",
          8070 => x"ca3f82b6",
          8071 => x"98085582",
          8072 => x"b698088c",
          8073 => x"387851ff",
          8074 => x"b5aa3f82",
          8075 => x"b6980855",
          8076 => x"7482b698",
          8077 => x"0ca83d0d",
          8078 => x"04ed3d0d",
          8079 => x"0280db05",
          8080 => x"33028405",
          8081 => x"80df0533",
          8082 => x"57578253",
          8083 => x"953dd005",
          8084 => x"52963d51",
          8085 => x"d2e93f82",
          8086 => x"b6980855",
          8087 => x"82b69808",
          8088 => x"80cf3878",
          8089 => x"5a655295",
          8090 => x"3dd40551",
          8091 => x"c9b53f82",
          8092 => x"b6980855",
          8093 => x"82b69808",
          8094 => x"b8380280",
          8095 => x"cf053381",
          8096 => x"a0065486",
          8097 => x"5573aa38",
          8098 => x"75a70661",
          8099 => x"71098b12",
          8100 => x"3371067a",
          8101 => x"74060751",
          8102 => x"57555674",
          8103 => x"8b153478",
          8104 => x"54810b83",
          8105 => x"15347851",
          8106 => x"ffb4a93f",
          8107 => x"82b69808",
          8108 => x"557482b6",
          8109 => x"980c953d",
          8110 => x"0d04ef3d",
          8111 => x"0d645682",
          8112 => x"53933dd0",
          8113 => x"0552943d",
          8114 => x"51d1f43f",
          8115 => x"82b69808",
          8116 => x"5582b698",
          8117 => x"0880cb38",
          8118 => x"76586352",
          8119 => x"933dd405",
          8120 => x"51c8c03f",
          8121 => x"82b69808",
          8122 => x"5582b698",
          8123 => x"08b43802",
          8124 => x"80c70533",
          8125 => x"81a00654",
          8126 => x"865573a6",
          8127 => x"38841622",
          8128 => x"86172271",
          8129 => x"902b0753",
          8130 => x"54961f51",
          8131 => x"ffb0c23f",
          8132 => x"7654810b",
          8133 => x"83153476",
          8134 => x"51ffb3b8",
          8135 => x"3f82b698",
          8136 => x"08557482",
          8137 => x"b6980c93",
          8138 => x"3d0d04ea",
          8139 => x"3d0d696b",
          8140 => x"5c5a8053",
          8141 => x"983dd005",
          8142 => x"52993d51",
          8143 => x"d1813f82",
          8144 => x"b6980882",
          8145 => x"b6980830",
          8146 => x"7082b698",
          8147 => x"08078025",
          8148 => x"51555779",
          8149 => x"802e8185",
          8150 => x"38817075",
          8151 => x"06555573",
          8152 => x"802e80f9",
          8153 => x"387b5d80",
          8154 => x"5f80528d",
          8155 => x"3d705254",
          8156 => x"ffbea93f",
          8157 => x"82b69808",
          8158 => x"5782b698",
          8159 => x"0880d138",
          8160 => x"74527351",
          8161 => x"c3dc3f82",
          8162 => x"b6980857",
          8163 => x"82b69808",
          8164 => x"bf3882b6",
          8165 => x"980882b6",
          8166 => x"9808655b",
          8167 => x"59567818",
          8168 => x"81197b18",
          8169 => x"56595574",
          8170 => x"33743481",
          8171 => x"16568a78",
          8172 => x"27ec388b",
          8173 => x"56751a54",
          8174 => x"80743475",
          8175 => x"802e9e38",
          8176 => x"ff16701b",
          8177 => x"70335155",
          8178 => x"5673a02e",
          8179 => x"e8388e39",
          8180 => x"76842e09",
          8181 => x"81068638",
          8182 => x"807a3480",
          8183 => x"57763070",
          8184 => x"78078025",
          8185 => x"51547a80",
          8186 => x"2e80c138",
          8187 => x"73802ebc",
          8188 => x"387ba011",
          8189 => x"085351ff",
          8190 => x"b1933f82",
          8191 => x"b6980857",
          8192 => x"82b69808",
          8193 => x"a7387b70",
          8194 => x"33555580",
          8195 => x"c3567383",
          8196 => x"2e8b3880",
          8197 => x"e4567384",
          8198 => x"2e8338a7",
          8199 => x"567515b4",
          8200 => x"0551ffad",
          8201 => x"e33f82b6",
          8202 => x"98087b0c",
          8203 => x"7682b698",
          8204 => x"0c983d0d",
          8205 => x"04e63d0d",
          8206 => x"82539c3d",
          8207 => x"ffb80552",
          8208 => x"9d3d51ce",
          8209 => x"fa3f82b6",
          8210 => x"980882b6",
          8211 => x"98085654",
          8212 => x"82b69808",
          8213 => x"8398388b",
          8214 => x"53a0528b",
          8215 => x"3d705259",
          8216 => x"ffaec03f",
          8217 => x"736d7033",
          8218 => x"7081ff06",
          8219 => x"52575557",
          8220 => x"9f742781",
          8221 => x"bc387858",
          8222 => x"7481ff06",
          8223 => x"6d81054e",
          8224 => x"705255ff",
          8225 => x"af893f82",
          8226 => x"b6980880",
          8227 => x"2ea5386c",
          8228 => x"70337053",
          8229 => x"5754ffae",
          8230 => x"fd3f82b6",
          8231 => x"9808802e",
          8232 => x"8d387488",
          8233 => x"2b76076d",
          8234 => x"81054e55",
          8235 => x"863982b6",
          8236 => x"980855ff",
          8237 => x"9f157083",
          8238 => x"ffff0651",
          8239 => x"54739926",
          8240 => x"8a38e015",
          8241 => x"7083ffff",
          8242 => x"06565480",
          8243 => x"ff752787",
          8244 => x"3882aee0",
          8245 => x"15335574",
          8246 => x"802ea338",
          8247 => x"745282b0",
          8248 => x"e051ffae",
          8249 => x"893f82b6",
          8250 => x"98089338",
          8251 => x"81ff7527",
          8252 => x"88387689",
          8253 => x"2688388b",
          8254 => x"398a7727",
          8255 => x"86388655",
          8256 => x"81ec3981",
          8257 => x"ff75278f",
          8258 => x"3874882a",
          8259 => x"54737870",
          8260 => x"81055a34",
          8261 => x"81175774",
          8262 => x"78708105",
          8263 => x"5a348117",
          8264 => x"6d703370",
          8265 => x"81ff0652",
          8266 => x"57555773",
          8267 => x"9f26fec8",
          8268 => x"388b3d33",
          8269 => x"54865573",
          8270 => x"81e52e81",
          8271 => x"b1387680",
          8272 => x"2e993802",
          8273 => x"a7055576",
          8274 => x"15703351",
          8275 => x"5473a02e",
          8276 => x"09810687",
          8277 => x"38ff1757",
          8278 => x"76ed3879",
          8279 => x"41804380",
          8280 => x"52913d70",
          8281 => x"5255ffba",
          8282 => x"b33f82b6",
          8283 => x"98085482",
          8284 => x"b6980880",
          8285 => x"f7388152",
          8286 => x"7451ffbf",
          8287 => x"e53f82b6",
          8288 => x"98085482",
          8289 => x"b698088d",
          8290 => x"387680c4",
          8291 => x"386754e5",
          8292 => x"743480c6",
          8293 => x"3982b698",
          8294 => x"08842e09",
          8295 => x"810680cc",
          8296 => x"38805476",
          8297 => x"742e80c4",
          8298 => x"38815274",
          8299 => x"51ffbdb0",
          8300 => x"3f82b698",
          8301 => x"085482b6",
          8302 => x"9808b138",
          8303 => x"a05382b6",
          8304 => x"98085267",
          8305 => x"51ffabdb",
          8306 => x"3f675488",
          8307 => x"0b8b1534",
          8308 => x"8b537852",
          8309 => x"6751ffab",
          8310 => x"a73f7954",
          8311 => x"810b8315",
          8312 => x"347951ff",
          8313 => x"adee3f82",
          8314 => x"b6980854",
          8315 => x"73557482",
          8316 => x"b6980c9c",
          8317 => x"3d0d04f2",
          8318 => x"3d0d6062",
          8319 => x"02880580",
          8320 => x"cb053393",
          8321 => x"3dfc0555",
          8322 => x"7254405e",
          8323 => x"5ad2da3f",
          8324 => x"82b69808",
          8325 => x"5882b698",
          8326 => x"0882bd38",
          8327 => x"911a3358",
          8328 => x"7782b538",
          8329 => x"7c802e97",
          8330 => x"388c1a08",
          8331 => x"59789038",
          8332 => x"901a3370",
          8333 => x"812a7081",
          8334 => x"06515555",
          8335 => x"73903887",
          8336 => x"54829739",
          8337 => x"82588290",
          8338 => x"39815882",
          8339 => x"8b397e8a",
          8340 => x"11227089",
          8341 => x"2b70557f",
          8342 => x"54565656",
          8343 => x"fec2a43f",
          8344 => x"ff147d06",
          8345 => x"70307072",
          8346 => x"079f2a82",
          8347 => x"b6980805",
          8348 => x"8c19087c",
          8349 => x"405a5d55",
          8350 => x"55817727",
          8351 => x"88389816",
          8352 => x"08772683",
          8353 => x"38825776",
          8354 => x"77565980",
          8355 => x"56745279",
          8356 => x"51ffae99",
          8357 => x"3f81157f",
          8358 => x"55559814",
          8359 => x"08752683",
          8360 => x"38825582",
          8361 => x"b6980881",
          8362 => x"2eff9938",
          8363 => x"82b69808",
          8364 => x"ff2eff95",
          8365 => x"3882b698",
          8366 => x"088e3881",
          8367 => x"1656757b",
          8368 => x"2e098106",
          8369 => x"87389339",
          8370 => x"74598056",
          8371 => x"74772e09",
          8372 => x"8106ffb9",
          8373 => x"38875880",
          8374 => x"ff397d80",
          8375 => x"2eba3878",
          8376 => x"7b55557a",
          8377 => x"802eb438",
          8378 => x"81155673",
          8379 => x"812e0981",
          8380 => x"068338ff",
          8381 => x"56755374",
          8382 => x"527e51ff",
          8383 => x"afa83f82",
          8384 => x"b6980858",
          8385 => x"82b69808",
          8386 => x"80ce3874",
          8387 => x"8116ff16",
          8388 => x"56565c73",
          8389 => x"d3388439",
          8390 => x"ff195c7e",
          8391 => x"7c8c120c",
          8392 => x"557d802e",
          8393 => x"b3387888",
          8394 => x"1b0c7c8c",
          8395 => x"1b0c901a",
          8396 => x"3380c007",
          8397 => x"5473901b",
          8398 => x"34981508",
          8399 => x"fe059016",
          8400 => x"08575475",
          8401 => x"74269138",
          8402 => x"757b3190",
          8403 => x"160c8415",
          8404 => x"33810754",
          8405 => x"73841634",
          8406 => x"77547382",
          8407 => x"b6980c90",
          8408 => x"3d0d04e9",
          8409 => x"3d0d6b6d",
          8410 => x"02880580",
          8411 => x"eb05339d",
          8412 => x"3d545a5c",
          8413 => x"59c5bd3f",
          8414 => x"8b56800b",
          8415 => x"82b69808",
          8416 => x"248bf838",
          8417 => x"82b69808",
          8418 => x"842982cd",
          8419 => x"d0057008",
          8420 => x"51557480",
          8421 => x"2e843880",
          8422 => x"753482b6",
          8423 => x"980881ff",
          8424 => x"065f8152",
          8425 => x"7e51ffa0",
          8426 => x"d03f82b6",
          8427 => x"980881ff",
          8428 => x"06708106",
          8429 => x"56578356",
          8430 => x"748bc038",
          8431 => x"76822a70",
          8432 => x"81065155",
          8433 => x"8a56748b",
          8434 => x"b238993d",
          8435 => x"fc055383",
          8436 => x"527e51ff",
          8437 => x"a4f03f82",
          8438 => x"b6980899",
          8439 => x"38675574",
          8440 => x"802e9238",
          8441 => x"74828080",
          8442 => x"268b38ff",
          8443 => x"15750655",
          8444 => x"74802e83",
          8445 => x"38814878",
          8446 => x"802e8738",
          8447 => x"84807926",
          8448 => x"92387881",
          8449 => x"800a268b",
          8450 => x"38ff1979",
          8451 => x"06557480",
          8452 => x"2e863893",
          8453 => x"568ae439",
          8454 => x"78892a6e",
          8455 => x"892a7089",
          8456 => x"2b775948",
          8457 => x"43597a83",
          8458 => x"38815661",
          8459 => x"30708025",
          8460 => x"77075155",
          8461 => x"9156748a",
          8462 => x"c238993d",
          8463 => x"f8055381",
          8464 => x"527e51ff",
          8465 => x"a4803f81",
          8466 => x"5682b698",
          8467 => x"088aac38",
          8468 => x"77832a70",
          8469 => x"770682b6",
          8470 => x"98084356",
          8471 => x"45748338",
          8472 => x"bf416655",
          8473 => x"8e566075",
          8474 => x"268a9038",
          8475 => x"74613170",
          8476 => x"485580ff",
          8477 => x"75278a83",
          8478 => x"38935678",
          8479 => x"81802689",
          8480 => x"fa387781",
          8481 => x"2a708106",
          8482 => x"56437480",
          8483 => x"2e953877",
          8484 => x"87065574",
          8485 => x"822e838d",
          8486 => x"38778106",
          8487 => x"5574802e",
          8488 => x"83833877",
          8489 => x"81065593",
          8490 => x"56825e74",
          8491 => x"802e89cb",
          8492 => x"38785a7d",
          8493 => x"832e0981",
          8494 => x"0680e138",
          8495 => x"78ae3866",
          8496 => x"912a5781",
          8497 => x"0b82b184",
          8498 => x"22565a74",
          8499 => x"802e9d38",
          8500 => x"74772698",
          8501 => x"3882b184",
          8502 => x"56791082",
          8503 => x"17702257",
          8504 => x"575a7480",
          8505 => x"2e863876",
          8506 => x"7527ee38",
          8507 => x"79526651",
          8508 => x"febd903f",
          8509 => x"82b69808",
          8510 => x"84298487",
          8511 => x"0570892a",
          8512 => x"5e55a05c",
          8513 => x"800b82b6",
          8514 => x"9808fc80",
          8515 => x"8a055644",
          8516 => x"fdfff00a",
          8517 => x"752780ec",
          8518 => x"3888d339",
          8519 => x"78ae3866",
          8520 => x"8c2a5781",
          8521 => x"0b82b0f4",
          8522 => x"22565a74",
          8523 => x"802e9d38",
          8524 => x"74772698",
          8525 => x"3882b0f4",
          8526 => x"56791082",
          8527 => x"17702257",
          8528 => x"575a7480",
          8529 => x"2e863876",
          8530 => x"7527ee38",
          8531 => x"79526651",
          8532 => x"febcb03f",
          8533 => x"82b69808",
          8534 => x"10840557",
          8535 => x"82b69808",
          8536 => x"9ff52696",
          8537 => x"38810b82",
          8538 => x"b6980810",
          8539 => x"82b69808",
          8540 => x"05711172",
          8541 => x"2a830559",
          8542 => x"565e83ff",
          8543 => x"17892a5d",
          8544 => x"815ca044",
          8545 => x"601c7d11",
          8546 => x"65056970",
          8547 => x"12ff0571",
          8548 => x"30707206",
          8549 => x"74315c52",
          8550 => x"59575940",
          8551 => x"7d832e09",
          8552 => x"81068938",
          8553 => x"761c6018",
          8554 => x"415c8439",
          8555 => x"761d5d79",
          8556 => x"90291870",
          8557 => x"62316858",
          8558 => x"51557476",
          8559 => x"2687af38",
          8560 => x"757c317d",
          8561 => x"317a5370",
          8562 => x"65315255",
          8563 => x"febbb43f",
          8564 => x"82b69808",
          8565 => x"587d832e",
          8566 => x"0981069b",
          8567 => x"3882b698",
          8568 => x"0883fff5",
          8569 => x"2680dd38",
          8570 => x"78878338",
          8571 => x"79812a59",
          8572 => x"78fdbe38",
          8573 => x"86f8397d",
          8574 => x"822e0981",
          8575 => x"0680c538",
          8576 => x"83fff50b",
          8577 => x"82b69808",
          8578 => x"27a03878",
          8579 => x"8f38791a",
          8580 => x"557480c0",
          8581 => x"26863874",
          8582 => x"59fd9639",
          8583 => x"62810655",
          8584 => x"74802e8f",
          8585 => x"38835efd",
          8586 => x"883982b6",
          8587 => x"98089ff5",
          8588 => x"26923878",
          8589 => x"86b83879",
          8590 => x"1a598180",
          8591 => x"7927fcf1",
          8592 => x"3886ab39",
          8593 => x"80557d81",
          8594 => x"2e098106",
          8595 => x"83387d55",
          8596 => x"9ff57827",
          8597 => x"8b387481",
          8598 => x"06558e56",
          8599 => x"74869c38",
          8600 => x"84805380",
          8601 => x"527a51ff",
          8602 => x"a2b93f8b",
          8603 => x"5382af9c",
          8604 => x"527a51ff",
          8605 => x"a28a3f84",
          8606 => x"80528b1b",
          8607 => x"51ffa1b3",
          8608 => x"3f798d1c",
          8609 => x"347b83ff",
          8610 => x"ff06528e",
          8611 => x"1b51ffa1",
          8612 => x"a23f810b",
          8613 => x"901c347d",
          8614 => x"83327030",
          8615 => x"70962a84",
          8616 => x"80065451",
          8617 => x"55911b51",
          8618 => x"ffa1883f",
          8619 => x"66557483",
          8620 => x"ffff2690",
          8621 => x"387483ff",
          8622 => x"ff065293",
          8623 => x"1b51ffa0",
          8624 => x"f23f8a39",
          8625 => x"7452a01b",
          8626 => x"51ffa185",
          8627 => x"3ff80b95",
          8628 => x"1c34bf52",
          8629 => x"981b51ff",
          8630 => x"a0d93f81",
          8631 => x"ff529a1b",
          8632 => x"51ffa0cf",
          8633 => x"3f60529c",
          8634 => x"1b51ffa0",
          8635 => x"e43f7d83",
          8636 => x"2e098106",
          8637 => x"80cb3882",
          8638 => x"88b20a52",
          8639 => x"80c31b51",
          8640 => x"ffa0ce3f",
          8641 => x"7c52a41b",
          8642 => x"51ffa0c5",
          8643 => x"3f8252ac",
          8644 => x"1b51ffa0",
          8645 => x"bc3f8152",
          8646 => x"b01b51ff",
          8647 => x"a0953f86",
          8648 => x"52b21b51",
          8649 => x"ffa08c3f",
          8650 => x"ff800b80",
          8651 => x"c01c34a9",
          8652 => x"0b80c21c",
          8653 => x"34935382",
          8654 => x"afa85280",
          8655 => x"c71b51ae",
          8656 => x"398288b2",
          8657 => x"0a52a71b",
          8658 => x"51ffa085",
          8659 => x"3f7c83ff",
          8660 => x"ff065296",
          8661 => x"1b51ff9f",
          8662 => x"da3fff80",
          8663 => x"0ba41c34",
          8664 => x"a90ba61c",
          8665 => x"34935382",
          8666 => x"afbc52ab",
          8667 => x"1b51ffa0",
          8668 => x"8f3f82d4",
          8669 => x"d55283fe",
          8670 => x"1b705259",
          8671 => x"ff9fb43f",
          8672 => x"81546053",
          8673 => x"7a527e51",
          8674 => x"ff9bd73f",
          8675 => x"815682b6",
          8676 => x"980883e7",
          8677 => x"387d832e",
          8678 => x"09810680",
          8679 => x"ee387554",
          8680 => x"60860553",
          8681 => x"7a527e51",
          8682 => x"ff9bb73f",
          8683 => x"84805380",
          8684 => x"527a51ff",
          8685 => x"9fed3f84",
          8686 => x"8b85a4d2",
          8687 => x"527a51ff",
          8688 => x"9f8f3f86",
          8689 => x"8a85e4f2",
          8690 => x"5283e41b",
          8691 => x"51ff9f81",
          8692 => x"3fff1852",
          8693 => x"83e81b51",
          8694 => x"ff9ef63f",
          8695 => x"825283ec",
          8696 => x"1b51ff9e",
          8697 => x"ec3f82d4",
          8698 => x"d5527851",
          8699 => x"ff9ec43f",
          8700 => x"75546087",
          8701 => x"05537a52",
          8702 => x"7e51ff9a",
          8703 => x"e53f7554",
          8704 => x"6016537a",
          8705 => x"527e51ff",
          8706 => x"9ad83f65",
          8707 => x"5380527a",
          8708 => x"51ff9f8f",
          8709 => x"3f7f5680",
          8710 => x"587d832e",
          8711 => x"0981069a",
          8712 => x"38f8527a",
          8713 => x"51ff9ea9",
          8714 => x"3fff5284",
          8715 => x"1b51ff9e",
          8716 => x"a03ff00a",
          8717 => x"52881b51",
          8718 => x"913987ff",
          8719 => x"fff8557d",
          8720 => x"812e8338",
          8721 => x"f8557452",
          8722 => x"7a51ff9e",
          8723 => x"843f7c55",
          8724 => x"61577462",
          8725 => x"26833874",
          8726 => x"57765475",
          8727 => x"537a527e",
          8728 => x"51ff99fe",
          8729 => x"3f82b698",
          8730 => x"08828738",
          8731 => x"84805382",
          8732 => x"b6980852",
          8733 => x"7a51ff9e",
          8734 => x"aa3f7616",
          8735 => x"75783156",
          8736 => x"5674cd38",
          8737 => x"81185877",
          8738 => x"802eff8d",
          8739 => x"3879557d",
          8740 => x"832e8338",
          8741 => x"63556157",
          8742 => x"74622683",
          8743 => x"38745776",
          8744 => x"5475537a",
          8745 => x"527e51ff",
          8746 => x"99b83f82",
          8747 => x"b6980881",
          8748 => x"c1387616",
          8749 => x"75783156",
          8750 => x"5674db38",
          8751 => x"8c567d83",
          8752 => x"2e933886",
          8753 => x"566683ff",
          8754 => x"ff268a38",
          8755 => x"84567d82",
          8756 => x"2e833881",
          8757 => x"56648106",
          8758 => x"587780fe",
          8759 => x"38848053",
          8760 => x"77527a51",
          8761 => x"ff9dbc3f",
          8762 => x"82d4d552",
          8763 => x"7851ff9c",
          8764 => x"c23f83be",
          8765 => x"1b557775",
          8766 => x"34810b81",
          8767 => x"1634810b",
          8768 => x"82163477",
          8769 => x"83163475",
          8770 => x"84163460",
          8771 => x"67055680",
          8772 => x"fdc15275",
          8773 => x"51feb4eb",
          8774 => x"3ffe0b85",
          8775 => x"163482b6",
          8776 => x"9808822a",
          8777 => x"bf075675",
          8778 => x"86163482",
          8779 => x"b6980887",
          8780 => x"16346052",
          8781 => x"83c61b51",
          8782 => x"ff9c963f",
          8783 => x"665283ca",
          8784 => x"1b51ff9c",
          8785 => x"8c3f8154",
          8786 => x"77537a52",
          8787 => x"7e51ff98",
          8788 => x"913f8156",
          8789 => x"82b69808",
          8790 => x"a2388053",
          8791 => x"80527e51",
          8792 => x"ff99e33f",
          8793 => x"815682b6",
          8794 => x"98089038",
          8795 => x"89398e56",
          8796 => x"8a398156",
          8797 => x"863982b6",
          8798 => x"98085675",
          8799 => x"82b6980c",
          8800 => x"993d0d04",
          8801 => x"f53d0d7d",
          8802 => x"605b5980",
          8803 => x"7960ff05",
          8804 => x"5a575776",
          8805 => x"7825b438",
          8806 => x"8d3df811",
          8807 => x"55558153",
          8808 => x"fc155279",
          8809 => x"51c9dc3f",
          8810 => x"7a812e09",
          8811 => x"81069c38",
          8812 => x"8c3d3355",
          8813 => x"748d2edb",
          8814 => x"38747670",
          8815 => x"81055834",
          8816 => x"81175774",
          8817 => x"8a2e0981",
          8818 => x"06c93880",
          8819 => x"76347855",
          8820 => x"76833876",
          8821 => x"557482b6",
          8822 => x"980c8d3d",
          8823 => x"0d04f73d",
          8824 => x"0d7b0284",
          8825 => x"05b30533",
          8826 => x"5957778a",
          8827 => x"2e098106",
          8828 => x"87388d52",
          8829 => x"7651e73f",
          8830 => x"84170856",
          8831 => x"807624be",
          8832 => x"38881708",
          8833 => x"77178c05",
          8834 => x"56597775",
          8835 => x"34811656",
          8836 => x"bb7625a1",
          8837 => x"388b3dfc",
          8838 => x"05547553",
          8839 => x"8c175276",
          8840 => x"0851cbdc",
          8841 => x"3f797632",
          8842 => x"70307072",
          8843 => x"079f2a70",
          8844 => x"30535156",
          8845 => x"56758418",
          8846 => x"0c811988",
          8847 => x"180c8b3d",
          8848 => x"0d04f93d",
          8849 => x"0d798411",
          8850 => x"08565680",
          8851 => x"7524a738",
          8852 => x"893dfc05",
          8853 => x"5474538c",
          8854 => x"16527508",
          8855 => x"51cba13f",
          8856 => x"82b69808",
          8857 => x"91388416",
          8858 => x"08782e09",
          8859 => x"81068738",
          8860 => x"88160855",
          8861 => x"8339ff55",
          8862 => x"7482b698",
          8863 => x"0c893d0d",
          8864 => x"04fd3d0d",
          8865 => x"755480cc",
          8866 => x"53805273",
          8867 => x"51ff9a93",
          8868 => x"3f76740c",
          8869 => x"853d0d04",
          8870 => x"ea3d0d02",
          8871 => x"80e30533",
          8872 => x"6a53863d",
          8873 => x"70535454",
          8874 => x"d83f7352",
          8875 => x"7251feae",
          8876 => x"3f7251ff",
          8877 => x"8d3f983d",
          8878 => x"0d040000",
          8879 => x"00ffffff",
          8880 => x"ff00ffff",
          8881 => x"ffff00ff",
          8882 => x"ffffff00",
          8883 => x"00002baa",
          8884 => x"00002b2e",
          8885 => x"00002b35",
          8886 => x"00002b3c",
          8887 => x"00002b43",
          8888 => x"00002b4a",
          8889 => x"00002b51",
          8890 => x"00002b58",
          8891 => x"00002b5f",
          8892 => x"00002b66",
          8893 => x"00002b6d",
          8894 => x"00002b74",
          8895 => x"00002b7a",
          8896 => x"00002b80",
          8897 => x"00002b86",
          8898 => x"00002b8c",
          8899 => x"00002b92",
          8900 => x"00002b98",
          8901 => x"00002b9e",
          8902 => x"00002ba4",
          8903 => x"00004171",
          8904 => x"00004177",
          8905 => x"0000417d",
          8906 => x"00004183",
          8907 => x"00004189",
          8908 => x"00004767",
          8909 => x"00004867",
          8910 => x"00004978",
          8911 => x"00004bd0",
          8912 => x"0000484f",
          8913 => x"0000463c",
          8914 => x"00004a40",
          8915 => x"00004ba1",
          8916 => x"00004a83",
          8917 => x"00004b19",
          8918 => x"00004a9f",
          8919 => x"00004922",
          8920 => x"0000463c",
          8921 => x"00004978",
          8922 => x"000049a1",
          8923 => x"00004a40",
          8924 => x"0000463c",
          8925 => x"0000463c",
          8926 => x"00004a9f",
          8927 => x"00004b19",
          8928 => x"00004ba1",
          8929 => x"00004bd0",
          8930 => x"00000e31",
          8931 => x"0000171a",
          8932 => x"0000171a",
          8933 => x"00000e60",
          8934 => x"0000171a",
          8935 => x"0000171a",
          8936 => x"0000171a",
          8937 => x"0000171a",
          8938 => x"0000171a",
          8939 => x"0000171a",
          8940 => x"0000171a",
          8941 => x"00000e1d",
          8942 => x"0000171a",
          8943 => x"00000e48",
          8944 => x"00000e78",
          8945 => x"0000171a",
          8946 => x"0000171a",
          8947 => x"0000171a",
          8948 => x"0000171a",
          8949 => x"0000171a",
          8950 => x"0000171a",
          8951 => x"0000171a",
          8952 => x"0000171a",
          8953 => x"0000171a",
          8954 => x"0000171a",
          8955 => x"0000171a",
          8956 => x"0000171a",
          8957 => x"0000171a",
          8958 => x"0000171a",
          8959 => x"0000171a",
          8960 => x"0000171a",
          8961 => x"0000171a",
          8962 => x"0000171a",
          8963 => x"0000171a",
          8964 => x"0000171a",
          8965 => x"0000171a",
          8966 => x"0000171a",
          8967 => x"0000171a",
          8968 => x"0000171a",
          8969 => x"0000171a",
          8970 => x"0000171a",
          8971 => x"0000171a",
          8972 => x"0000171a",
          8973 => x"0000171a",
          8974 => x"0000171a",
          8975 => x"0000171a",
          8976 => x"0000171a",
          8977 => x"0000171a",
          8978 => x"0000171a",
          8979 => x"0000171a",
          8980 => x"0000171a",
          8981 => x"00000fa8",
          8982 => x"0000171a",
          8983 => x"0000171a",
          8984 => x"0000171a",
          8985 => x"0000171a",
          8986 => x"00001116",
          8987 => x"0000171a",
          8988 => x"0000171a",
          8989 => x"0000171a",
          8990 => x"0000171a",
          8991 => x"0000171a",
          8992 => x"0000171a",
          8993 => x"0000171a",
          8994 => x"0000171a",
          8995 => x"0000171a",
          8996 => x"0000171a",
          8997 => x"00000ed8",
          8998 => x"0000103f",
          8999 => x"00000eaf",
          9000 => x"00000eaf",
          9001 => x"00000eaf",
          9002 => x"0000171a",
          9003 => x"0000103f",
          9004 => x"0000171a",
          9005 => x"0000171a",
          9006 => x"00000e98",
          9007 => x"0000171a",
          9008 => x"0000171a",
          9009 => x"000010ec",
          9010 => x"000010f7",
          9011 => x"0000171a",
          9012 => x"0000171a",
          9013 => x"00000f11",
          9014 => x"0000171a",
          9015 => x"0000111f",
          9016 => x"0000171a",
          9017 => x"0000171a",
          9018 => x"00001116",
          9019 => x"64696e69",
          9020 => x"74000000",
          9021 => x"64696f63",
          9022 => x"746c0000",
          9023 => x"66696e69",
          9024 => x"74000000",
          9025 => x"666c6f61",
          9026 => x"64000000",
          9027 => x"66657865",
          9028 => x"63000000",
          9029 => x"6d636c65",
          9030 => x"61720000",
          9031 => x"6d636f70",
          9032 => x"79000000",
          9033 => x"6d646966",
          9034 => x"66000000",
          9035 => x"6d64756d",
          9036 => x"70000000",
          9037 => x"6d656200",
          9038 => x"6d656800",
          9039 => x"6d657700",
          9040 => x"68696400",
          9041 => x"68696500",
          9042 => x"68666400",
          9043 => x"68666500",
          9044 => x"63616c6c",
          9045 => x"00000000",
          9046 => x"6a6d7000",
          9047 => x"72657374",
          9048 => x"61727400",
          9049 => x"72657365",
          9050 => x"74000000",
          9051 => x"696e666f",
          9052 => x"00000000",
          9053 => x"74657374",
          9054 => x"00000000",
          9055 => x"74626173",
          9056 => x"69630000",
          9057 => x"6d626173",
          9058 => x"69630000",
          9059 => x"6b696c6f",
          9060 => x"00000000",
          9061 => x"65640000",
          9062 => x"4469736b",
          9063 => x"20457272",
          9064 => x"6f720000",
          9065 => x"496e7465",
          9066 => x"726e616c",
          9067 => x"20657272",
          9068 => x"6f722e00",
          9069 => x"4469736b",
          9070 => x"206e6f74",
          9071 => x"20726561",
          9072 => x"64792e00",
          9073 => x"4e6f2066",
          9074 => x"696c6520",
          9075 => x"666f756e",
          9076 => x"642e0000",
          9077 => x"4e6f2070",
          9078 => x"61746820",
          9079 => x"666f756e",
          9080 => x"642e0000",
          9081 => x"496e7661",
          9082 => x"6c696420",
          9083 => x"66696c65",
          9084 => x"6e616d65",
          9085 => x"2e000000",
          9086 => x"41636365",
          9087 => x"73732064",
          9088 => x"656e6965",
          9089 => x"642e0000",
          9090 => x"46696c65",
          9091 => x"20616c72",
          9092 => x"65616479",
          9093 => x"20657869",
          9094 => x"7374732e",
          9095 => x"00000000",
          9096 => x"46696c65",
          9097 => x"2068616e",
          9098 => x"646c6520",
          9099 => x"696e7661",
          9100 => x"6c69642e",
          9101 => x"00000000",
          9102 => x"53442069",
          9103 => x"73207772",
          9104 => x"69746520",
          9105 => x"70726f74",
          9106 => x"65637465",
          9107 => x"642e0000",
          9108 => x"44726976",
          9109 => x"65206e75",
          9110 => x"6d626572",
          9111 => x"20697320",
          9112 => x"696e7661",
          9113 => x"6c69642e",
          9114 => x"00000000",
          9115 => x"4469736b",
          9116 => x"206e6f74",
          9117 => x"20656e61",
          9118 => x"626c6564",
          9119 => x"2e000000",
          9120 => x"4e6f2063",
          9121 => x"6f6d7061",
          9122 => x"7469626c",
          9123 => x"65206669",
          9124 => x"6c657379",
          9125 => x"7374656d",
          9126 => x"20666f75",
          9127 => x"6e64206f",
          9128 => x"6e206469",
          9129 => x"736b2e00",
          9130 => x"466f726d",
          9131 => x"61742061",
          9132 => x"626f7274",
          9133 => x"65642e00",
          9134 => x"54696d65",
          9135 => x"6f75742c",
          9136 => x"206f7065",
          9137 => x"72617469",
          9138 => x"6f6e2063",
          9139 => x"616e6365",
          9140 => x"6c6c6564",
          9141 => x"2e000000",
          9142 => x"46696c65",
          9143 => x"20697320",
          9144 => x"6c6f636b",
          9145 => x"65642e00",
          9146 => x"496e7375",
          9147 => x"66666963",
          9148 => x"69656e74",
          9149 => x"206d656d",
          9150 => x"6f72792e",
          9151 => x"00000000",
          9152 => x"546f6f20",
          9153 => x"6d616e79",
          9154 => x"206f7065",
          9155 => x"6e206669",
          9156 => x"6c65732e",
          9157 => x"00000000",
          9158 => x"50617261",
          9159 => x"6d657465",
          9160 => x"72732069",
          9161 => x"6e636f72",
          9162 => x"72656374",
          9163 => x"2e000000",
          9164 => x"53756363",
          9165 => x"6573732e",
          9166 => x"00000000",
          9167 => x"556e6b6e",
          9168 => x"6f776e20",
          9169 => x"6572726f",
          9170 => x"722e0000",
          9171 => x"0a256c75",
          9172 => x"20627974",
          9173 => x"65732025",
          9174 => x"73206174",
          9175 => x"20256c75",
          9176 => x"20627974",
          9177 => x"65732f73",
          9178 => x"65632e0a",
          9179 => x"00000000",
          9180 => x"72656164",
          9181 => x"00000000",
          9182 => x"303d2530",
          9183 => x"386c782c",
          9184 => x"20313d25",
          9185 => x"30386c78",
          9186 => x"2c20323d",
          9187 => x"2530386c",
          9188 => x"782c205f",
          9189 => x"494f423d",
          9190 => x"2530386c",
          9191 => x"78202530",
          9192 => x"386c7820",
          9193 => x"2530386c",
          9194 => x"780a0000",
          9195 => x"2530386c",
          9196 => x"58000000",
          9197 => x"3a202000",
          9198 => x"25303458",
          9199 => x"00000000",
          9200 => x"20202020",
          9201 => x"20202020",
          9202 => x"00000000",
          9203 => x"25303258",
          9204 => x"00000000",
          9205 => x"20200000",
          9206 => x"207c0000",
          9207 => x"7c000000",
          9208 => x"7a4f5300",
          9209 => x"0a2a2a20",
          9210 => x"25732028",
          9211 => x"00000000",
          9212 => x"30322f30",
          9213 => x"352f3230",
          9214 => x"32300000",
          9215 => x"76312e30",
          9216 => x"32000000",
          9217 => x"205a5055",
          9218 => x"2c207265",
          9219 => x"76202530",
          9220 => x"32782920",
          9221 => x"25732025",
          9222 => x"73202a2a",
          9223 => x"0a0a0000",
          9224 => x"5a505520",
          9225 => x"496e7465",
          9226 => x"72727570",
          9227 => x"74204861",
          9228 => x"6e646c65",
          9229 => x"72000000",
          9230 => x"54696d65",
          9231 => x"7220696e",
          9232 => x"74657272",
          9233 => x"75707400",
          9234 => x"50533220",
          9235 => x"696e7465",
          9236 => x"72727570",
          9237 => x"74000000",
          9238 => x"494f4354",
          9239 => x"4c205244",
          9240 => x"20696e74",
          9241 => x"65727275",
          9242 => x"70740000",
          9243 => x"494f4354",
          9244 => x"4c205752",
          9245 => x"20696e74",
          9246 => x"65727275",
          9247 => x"70740000",
          9248 => x"55415254",
          9249 => x"30205258",
          9250 => x"20696e74",
          9251 => x"65727275",
          9252 => x"70740000",
          9253 => x"55415254",
          9254 => x"30205458",
          9255 => x"20696e74",
          9256 => x"65727275",
          9257 => x"70740000",
          9258 => x"55415254",
          9259 => x"31205258",
          9260 => x"20696e74",
          9261 => x"65727275",
          9262 => x"70740000",
          9263 => x"55415254",
          9264 => x"31205458",
          9265 => x"20696e74",
          9266 => x"65727275",
          9267 => x"70740000",
          9268 => x"53657474",
          9269 => x"696e6720",
          9270 => x"75702074",
          9271 => x"696d6572",
          9272 => x"2e2e2e00",
          9273 => x"456e6162",
          9274 => x"6c696e67",
          9275 => x"2074696d",
          9276 => x"65722e2e",
          9277 => x"2e000000",
          9278 => x"6175746f",
          9279 => x"65786563",
          9280 => x"2e626174",
          9281 => x"00000000",
          9282 => x"7a4f532e",
          9283 => x"68737400",
          9284 => x"303a0000",
          9285 => x"4661696c",
          9286 => x"65642074",
          9287 => x"6f20696e",
          9288 => x"69746961",
          9289 => x"6c697365",
          9290 => x"20736420",
          9291 => x"63617264",
          9292 => x"20302c20",
          9293 => x"706c6561",
          9294 => x"73652069",
          9295 => x"6e697420",
          9296 => x"6d616e75",
          9297 => x"616c6c79",
          9298 => x"2e000000",
          9299 => x"2a200000",
          9300 => x"436c6561",
          9301 => x"72696e67",
          9302 => x"2e2e2e2e",
          9303 => x"00000000",
          9304 => x"436f7079",
          9305 => x"696e672e",
          9306 => x"2e2e0000",
          9307 => x"436f6d70",
          9308 => x"6172696e",
          9309 => x"672e2e2e",
          9310 => x"00000000",
          9311 => x"2530386c",
          9312 => x"78282530",
          9313 => x"3878292d",
          9314 => x"3e253038",
          9315 => x"6c782825",
          9316 => x"30387829",
          9317 => x"0a000000",
          9318 => x"44756d70",
          9319 => x"204d656d",
          9320 => x"6f727900",
          9321 => x"0a436f6d",
          9322 => x"706c6574",
          9323 => x"652e0000",
          9324 => x"2530386c",
          9325 => x"58202530",
          9326 => x"32582d00",
          9327 => x"3f3f3f00",
          9328 => x"2530386c",
          9329 => x"58202530",
          9330 => x"34582d00",
          9331 => x"2530386c",
          9332 => x"58202530",
          9333 => x"386c582d",
          9334 => x"00000000",
          9335 => x"45786563",
          9336 => x"7574696e",
          9337 => x"6720636f",
          9338 => x"64652040",
          9339 => x"20253038",
          9340 => x"6c78202e",
          9341 => x"2e2e0a00",
          9342 => x"43616c6c",
          9343 => x"696e6720",
          9344 => x"636f6465",
          9345 => x"20402025",
          9346 => x"30386c78",
          9347 => x"202e2e2e",
          9348 => x"0a000000",
          9349 => x"43616c6c",
          9350 => x"20726574",
          9351 => x"75726e65",
          9352 => x"6420636f",
          9353 => x"64652028",
          9354 => x"2564292e",
          9355 => x"0a000000",
          9356 => x"52657374",
          9357 => x"61727469",
          9358 => x"6e672061",
          9359 => x"70706c69",
          9360 => x"63617469",
          9361 => x"6f6e2e2e",
          9362 => x"2e000000",
          9363 => x"436f6c64",
          9364 => x"20726562",
          9365 => x"6f6f7469",
          9366 => x"6e672e2e",
          9367 => x"2e000000",
          9368 => x"5a505500",
          9369 => x"62696e00",
          9370 => x"25643a5c",
          9371 => x"25735c25",
          9372 => x"732e2573",
          9373 => x"00000000",
          9374 => x"25643a5c",
          9375 => x"25735c25",
          9376 => x"73000000",
          9377 => x"25643a5c",
          9378 => x"25730000",
          9379 => x"42616420",
          9380 => x"636f6d6d",
          9381 => x"616e642e",
          9382 => x"00000000",
          9383 => x"52756e6e",
          9384 => x"696e672e",
          9385 => x"2e2e0000",
          9386 => x"456e6162",
          9387 => x"6c696e67",
          9388 => x"20696e74",
          9389 => x"65727275",
          9390 => x"7074732e",
          9391 => x"2e2e0000",
          9392 => x"25642f25",
          9393 => x"642f2564",
          9394 => x"2025643a",
          9395 => x"25643a25",
          9396 => x"642e2564",
          9397 => x"25640a00",
          9398 => x"536f4320",
          9399 => x"436f6e66",
          9400 => x"69677572",
          9401 => x"6174696f",
          9402 => x"6e000000",
          9403 => x"20286672",
          9404 => x"6f6d2053",
          9405 => x"6f432063",
          9406 => x"6f6e6669",
          9407 => x"67290000",
          9408 => x"3a0a4465",
          9409 => x"76696365",
          9410 => x"7320696d",
          9411 => x"706c656d",
          9412 => x"656e7465",
          9413 => x"643a0000",
          9414 => x"20202020",
          9415 => x"57422053",
          9416 => x"4452414d",
          9417 => x"20202825",
          9418 => x"3038583a",
          9419 => x"25303858",
          9420 => x"292e0a00",
          9421 => x"20202020",
          9422 => x"53445241",
          9423 => x"4d202020",
          9424 => x"20202825",
          9425 => x"3038583a",
          9426 => x"25303858",
          9427 => x"292e0a00",
          9428 => x"20202020",
          9429 => x"494e534e",
          9430 => x"20425241",
          9431 => x"4d202825",
          9432 => x"3038583a",
          9433 => x"25303858",
          9434 => x"292e0a00",
          9435 => x"20202020",
          9436 => x"4252414d",
          9437 => x"20202020",
          9438 => x"20202825",
          9439 => x"3038583a",
          9440 => x"25303858",
          9441 => x"292e0a00",
          9442 => x"20202020",
          9443 => x"52414d20",
          9444 => x"20202020",
          9445 => x"20202825",
          9446 => x"3038583a",
          9447 => x"25303858",
          9448 => x"292e0a00",
          9449 => x"20202020",
          9450 => x"53442043",
          9451 => x"41524420",
          9452 => x"20202844",
          9453 => x"65766963",
          9454 => x"6573203d",
          9455 => x"25303264",
          9456 => x"292e0a00",
          9457 => x"20202020",
          9458 => x"54494d45",
          9459 => x"52312020",
          9460 => x"20202854",
          9461 => x"696d6572",
          9462 => x"7320203d",
          9463 => x"25303264",
          9464 => x"292e0a00",
          9465 => x"20202020",
          9466 => x"494e5452",
          9467 => x"20435452",
          9468 => x"4c202843",
          9469 => x"68616e6e",
          9470 => x"656c733d",
          9471 => x"25303264",
          9472 => x"292e0a00",
          9473 => x"20202020",
          9474 => x"57495348",
          9475 => x"424f4e45",
          9476 => x"20425553",
          9477 => x"00000000",
          9478 => x"20202020",
          9479 => x"57422049",
          9480 => x"32430000",
          9481 => x"20202020",
          9482 => x"494f4354",
          9483 => x"4c000000",
          9484 => x"20202020",
          9485 => x"50533200",
          9486 => x"20202020",
          9487 => x"53504900",
          9488 => x"41646472",
          9489 => x"65737365",
          9490 => x"733a0000",
          9491 => x"20202020",
          9492 => x"43505520",
          9493 => x"52657365",
          9494 => x"74205665",
          9495 => x"63746f72",
          9496 => x"20416464",
          9497 => x"72657373",
          9498 => x"203d2025",
          9499 => x"3038580a",
          9500 => x"00000000",
          9501 => x"20202020",
          9502 => x"43505520",
          9503 => x"4d656d6f",
          9504 => x"72792053",
          9505 => x"74617274",
          9506 => x"20416464",
          9507 => x"72657373",
          9508 => x"203d2025",
          9509 => x"3038580a",
          9510 => x"00000000",
          9511 => x"20202020",
          9512 => x"53746163",
          9513 => x"6b205374",
          9514 => x"61727420",
          9515 => x"41646472",
          9516 => x"65737320",
          9517 => x"20202020",
          9518 => x"203d2025",
          9519 => x"3038580a",
          9520 => x"00000000",
          9521 => x"4d697363",
          9522 => x"3a000000",
          9523 => x"20202020",
          9524 => x"5a505520",
          9525 => x"49642020",
          9526 => x"20202020",
          9527 => x"20202020",
          9528 => x"20202020",
          9529 => x"20202020",
          9530 => x"203d2025",
          9531 => x"3034580a",
          9532 => x"00000000",
          9533 => x"20202020",
          9534 => x"53797374",
          9535 => x"656d2043",
          9536 => x"6c6f636b",
          9537 => x"20467265",
          9538 => x"71202020",
          9539 => x"20202020",
          9540 => x"203d2025",
          9541 => x"642e2530",
          9542 => x"34644d48",
          9543 => x"7a0a0000",
          9544 => x"20202020",
          9545 => x"53445241",
          9546 => x"4d20436c",
          9547 => x"6f636b20",
          9548 => x"46726571",
          9549 => x"20202020",
          9550 => x"20202020",
          9551 => x"203d2025",
          9552 => x"642e2530",
          9553 => x"34644d48",
          9554 => x"7a0a0000",
          9555 => x"20202020",
          9556 => x"57697368",
          9557 => x"626f6e65",
          9558 => x"20534452",
          9559 => x"414d2043",
          9560 => x"6c6f636b",
          9561 => x"20467265",
          9562 => x"713d2025",
          9563 => x"642e2530",
          9564 => x"34644d48",
          9565 => x"7a0a0000",
          9566 => x"536d616c",
          9567 => x"6c000000",
          9568 => x"4d656469",
          9569 => x"756d0000",
          9570 => x"466c6578",
          9571 => x"00000000",
          9572 => x"45564f00",
          9573 => x"45564f6d",
          9574 => x"00000000",
          9575 => x"556e6b6e",
          9576 => x"6f776e00",
          9577 => x"00009700",
          9578 => x"01000000",
          9579 => x"00000002",
          9580 => x"000096fc",
          9581 => x"01000000",
          9582 => x"00000003",
          9583 => x"000096f8",
          9584 => x"01000000",
          9585 => x"00000004",
          9586 => x"000096f4",
          9587 => x"01000000",
          9588 => x"00000005",
          9589 => x"000096f0",
          9590 => x"01000000",
          9591 => x"00000006",
          9592 => x"000096ec",
          9593 => x"01000000",
          9594 => x"00000007",
          9595 => x"000096e8",
          9596 => x"01000000",
          9597 => x"00000001",
          9598 => x"000096e4",
          9599 => x"01000000",
          9600 => x"00000008",
          9601 => x"000096e0",
          9602 => x"01000000",
          9603 => x"0000000b",
          9604 => x"000096dc",
          9605 => x"01000000",
          9606 => x"00000009",
          9607 => x"000096d8",
          9608 => x"01000000",
          9609 => x"0000000a",
          9610 => x"000096d4",
          9611 => x"04000000",
          9612 => x"0000000d",
          9613 => x"000096d0",
          9614 => x"04000000",
          9615 => x"0000000c",
          9616 => x"000096cc",
          9617 => x"04000000",
          9618 => x"0000000e",
          9619 => x"000096c8",
          9620 => x"03000000",
          9621 => x"0000000f",
          9622 => x"000096c4",
          9623 => x"04000000",
          9624 => x"0000000f",
          9625 => x"000096c0",
          9626 => x"04000000",
          9627 => x"00000010",
          9628 => x"000096bc",
          9629 => x"04000000",
          9630 => x"00000011",
          9631 => x"000096b8",
          9632 => x"03000000",
          9633 => x"00000012",
          9634 => x"000096b4",
          9635 => x"03000000",
          9636 => x"00000013",
          9637 => x"000096b0",
          9638 => x"03000000",
          9639 => x"00000014",
          9640 => x"000096ac",
          9641 => x"03000000",
          9642 => x"00000015",
          9643 => x"1b5b4400",
          9644 => x"1b5b4300",
          9645 => x"1b5b4200",
          9646 => x"1b5b4100",
          9647 => x"1b5b367e",
          9648 => x"1b5b357e",
          9649 => x"1b5b347e",
          9650 => x"1b304600",
          9651 => x"1b5b337e",
          9652 => x"1b5b327e",
          9653 => x"1b5b317e",
          9654 => x"10000000",
          9655 => x"0e000000",
          9656 => x"0d000000",
          9657 => x"0b000000",
          9658 => x"08000000",
          9659 => x"06000000",
          9660 => x"05000000",
          9661 => x"04000000",
          9662 => x"03000000",
          9663 => x"02000000",
          9664 => x"01000000",
          9665 => x"68697374",
          9666 => x"6f727900",
          9667 => x"68697374",
          9668 => x"00000000",
          9669 => x"21000000",
          9670 => x"2530346c",
          9671 => x"75202025",
          9672 => x"730a0000",
          9673 => x"4661696c",
          9674 => x"65642074",
          9675 => x"6f207265",
          9676 => x"73657420",
          9677 => x"74686520",
          9678 => x"68697374",
          9679 => x"6f727920",
          9680 => x"66696c65",
          9681 => x"20746f20",
          9682 => x"454f462e",
          9683 => x"00000000",
          9684 => x"43616e6e",
          9685 => x"6f74206f",
          9686 => x"70656e2f",
          9687 => x"63726561",
          9688 => x"74652068",
          9689 => x"6973746f",
          9690 => x"72792066",
          9691 => x"696c652c",
          9692 => x"20646973",
          9693 => x"61626c69",
          9694 => x"6e672e00",
          9695 => x"53440000",
          9696 => x"222a2b2c",
          9697 => x"3a3b3c3d",
          9698 => x"3e3f5b5d",
          9699 => x"7c7f0000",
          9700 => x"46415400",
          9701 => x"46415433",
          9702 => x"32000000",
          9703 => x"ebfe904d",
          9704 => x"53444f53",
          9705 => x"352e3000",
          9706 => x"4e4f204e",
          9707 => x"414d4520",
          9708 => x"20202046",
          9709 => x"41543332",
          9710 => x"20202000",
          9711 => x"4e4f204e",
          9712 => x"414d4520",
          9713 => x"20202046",
          9714 => x"41542020",
          9715 => x"20202000",
          9716 => x"0000977c",
          9717 => x"00000000",
          9718 => x"00000000",
          9719 => x"00000000",
          9720 => x"809a4541",
          9721 => x"8e418f80",
          9722 => x"45454549",
          9723 => x"49498e8f",
          9724 => x"9092924f",
          9725 => x"994f5555",
          9726 => x"59999a9b",
          9727 => x"9c9d9e9f",
          9728 => x"41494f55",
          9729 => x"a5a5a6a7",
          9730 => x"a8a9aaab",
          9731 => x"acadaeaf",
          9732 => x"b0b1b2b3",
          9733 => x"b4b5b6b7",
          9734 => x"b8b9babb",
          9735 => x"bcbdbebf",
          9736 => x"c0c1c2c3",
          9737 => x"c4c5c6c7",
          9738 => x"c8c9cacb",
          9739 => x"cccdcecf",
          9740 => x"d0d1d2d3",
          9741 => x"d4d5d6d7",
          9742 => x"d8d9dadb",
          9743 => x"dcdddedf",
          9744 => x"e0e1e2e3",
          9745 => x"e4e5e6e7",
          9746 => x"e8e9eaeb",
          9747 => x"ecedeeef",
          9748 => x"f0f1f2f3",
          9749 => x"f4f5f6f7",
          9750 => x"f8f9fafb",
          9751 => x"fcfdfeff",
          9752 => x"2b2e2c3b",
          9753 => x"3d5b5d2f",
          9754 => x"5c222a3a",
          9755 => x"3c3e3f7c",
          9756 => x"7f000000",
          9757 => x"00010004",
          9758 => x"00100040",
          9759 => x"01000200",
          9760 => x"00000000",
          9761 => x"00010002",
          9762 => x"00040008",
          9763 => x"00100020",
          9764 => x"00000000",
          9765 => x"00000000",
          9766 => x"00008cec",
          9767 => x"01020100",
          9768 => x"00000000",
          9769 => x"00000000",
          9770 => x"00008cf4",
          9771 => x"01040100",
          9772 => x"00000000",
          9773 => x"00000000",
          9774 => x"00008cfc",
          9775 => x"01140300",
          9776 => x"00000000",
          9777 => x"00000000",
          9778 => x"00008d04",
          9779 => x"012b0300",
          9780 => x"00000000",
          9781 => x"00000000",
          9782 => x"00008d0c",
          9783 => x"01300300",
          9784 => x"00000000",
          9785 => x"00000000",
          9786 => x"00008d14",
          9787 => x"013c0400",
          9788 => x"00000000",
          9789 => x"00000000",
          9790 => x"00008d1c",
          9791 => x"013d0400",
          9792 => x"00000000",
          9793 => x"00000000",
          9794 => x"00008d24",
          9795 => x"013f0400",
          9796 => x"00000000",
          9797 => x"00000000",
          9798 => x"00008d2c",
          9799 => x"01400400",
          9800 => x"00000000",
          9801 => x"00000000",
          9802 => x"00008d34",
          9803 => x"01410400",
          9804 => x"00000000",
          9805 => x"00000000",
          9806 => x"00008d38",
          9807 => x"01420400",
          9808 => x"00000000",
          9809 => x"00000000",
          9810 => x"00008d3c",
          9811 => x"01430400",
          9812 => x"00000000",
          9813 => x"00000000",
          9814 => x"00008d40",
          9815 => x"01500500",
          9816 => x"00000000",
          9817 => x"00000000",
          9818 => x"00008d44",
          9819 => x"01510500",
          9820 => x"00000000",
          9821 => x"00000000",
          9822 => x"00008d48",
          9823 => x"01540500",
          9824 => x"00000000",
          9825 => x"00000000",
          9826 => x"00008d4c",
          9827 => x"01550500",
          9828 => x"00000000",
          9829 => x"00000000",
          9830 => x"00008d50",
          9831 => x"01790700",
          9832 => x"00000000",
          9833 => x"00000000",
          9834 => x"00008d58",
          9835 => x"01780700",
          9836 => x"00000000",
          9837 => x"00000000",
          9838 => x"00008d5c",
          9839 => x"01820800",
          9840 => x"00000000",
          9841 => x"00000000",
          9842 => x"00008d64",
          9843 => x"01830800",
          9844 => x"00000000",
          9845 => x"00000000",
          9846 => x"00008d6c",
          9847 => x"01850800",
          9848 => x"00000000",
          9849 => x"00000000",
          9850 => x"00008d74",
          9851 => x"01870800",
          9852 => x"00000000",
          9853 => x"00000000",
          9854 => x"00008d7c",
          9855 => x"018c0900",
          9856 => x"00000000",
          9857 => x"00000000",
          9858 => x"00008d84",
          9859 => x"018d0900",
          9860 => x"00000000",
          9861 => x"00000000",
          9862 => x"00008d8c",
          9863 => x"018e0900",
          9864 => x"00000000",
          9865 => x"00000000",
          9866 => x"00008d94",
          9867 => x"018f0900",
          9868 => x"00000000",
          9869 => x"00000000",
          9870 => x"00000000",
          9871 => x"00000000",
          9872 => x"00007fff",
          9873 => x"00000000",
          9874 => x"00007fff",
          9875 => x"00010000",
          9876 => x"00007fff",
          9877 => x"00010000",
          9878 => x"00810000",
          9879 => x"01000000",
          9880 => x"017fffff",
          9881 => x"00000000",
          9882 => x"00000000",
          9883 => x"00007800",
          9884 => x"00000000",
          9885 => x"05f5e100",
          9886 => x"05f5e100",
          9887 => x"05f5e100",
          9888 => x"00000000",
          9889 => x"01010101",
          9890 => x"01010101",
          9891 => x"01011001",
          9892 => x"01000000",
          9893 => x"00000000",
          9894 => x"00000000",
          9895 => x"00000000",
          9896 => x"00000000",
          9897 => x"00000000",
          9898 => x"00000000",
          9899 => x"00000000",
          9900 => x"00000000",
          9901 => x"00000000",
          9902 => x"00000000",
          9903 => x"00000000",
          9904 => x"00000000",
          9905 => x"00000000",
          9906 => x"00000000",
          9907 => x"00000000",
          9908 => x"00000000",
          9909 => x"00000000",
          9910 => x"00000000",
          9911 => x"00000000",
          9912 => x"00000000",
          9913 => x"00000000",
          9914 => x"00000000",
          9915 => x"00000000",
          9916 => x"00000000",
          9917 => x"00009704",
          9918 => x"01000000",
          9919 => x"0000970c",
          9920 => x"01000000",
          9921 => x"00009714",
          9922 => x"02000000",
          9923 => x"00000000",
          9924 => x"00000000",
          9925 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

