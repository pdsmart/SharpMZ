-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"ff",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"80",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"95",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"c3",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"c5",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"a4",
           386 => x"fe",
           387 => x"a4",
           388 => x"90",
           389 => x"a4",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"82",
           395 => x"82",
           396 => x"82",
           397 => x"af",
           398 => x"b6",
           399 => x"d0",
           400 => x"b6",
           401 => x"ad",
           402 => x"a4",
           403 => x"90",
           404 => x"a4",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"82",
           418 => x"82",
           419 => x"82",
           420 => x"96",
           421 => x"b6",
           422 => x"d0",
           423 => x"b6",
           424 => x"cd",
           425 => x"a4",
           426 => x"90",
           427 => x"a4",
           428 => x"a8",
           429 => x"a4",
           430 => x"90",
           431 => x"a4",
           432 => x"86",
           433 => x"a4",
           434 => x"90",
           435 => x"a4",
           436 => x"c3",
           437 => x"a4",
           438 => x"90",
           439 => x"a4",
           440 => x"ba",
           441 => x"a4",
           442 => x"90",
           443 => x"a4",
           444 => x"ed",
           445 => x"a4",
           446 => x"90",
           447 => x"a4",
           448 => x"9e",
           449 => x"a4",
           450 => x"90",
           451 => x"a4",
           452 => x"8f",
           453 => x"a4",
           454 => x"90",
           455 => x"a4",
           456 => x"83",
           457 => x"a4",
           458 => x"90",
           459 => x"a4",
           460 => x"80",
           461 => x"a4",
           462 => x"90",
           463 => x"a4",
           464 => x"9e",
           465 => x"a4",
           466 => x"90",
           467 => x"a4",
           468 => x"fe",
           469 => x"a4",
           470 => x"90",
           471 => x"a4",
           472 => x"f1",
           473 => x"a4",
           474 => x"90",
           475 => x"a4",
           476 => x"bd",
           477 => x"a4",
           478 => x"90",
           479 => x"a4",
           480 => x"dc",
           481 => x"a4",
           482 => x"90",
           483 => x"a4",
           484 => x"fb",
           485 => x"a4",
           486 => x"90",
           487 => x"a4",
           488 => x"e5",
           489 => x"a4",
           490 => x"90",
           491 => x"a4",
           492 => x"cb",
           493 => x"a4",
           494 => x"90",
           495 => x"a4",
           496 => x"b9",
           497 => x"a4",
           498 => x"90",
           499 => x"a4",
           500 => x"ff",
           501 => x"a4",
           502 => x"90",
           503 => x"a4",
           504 => x"b9",
           505 => x"a4",
           506 => x"90",
           507 => x"a4",
           508 => x"ba",
           509 => x"a4",
           510 => x"90",
           511 => x"a4",
           512 => x"ef",
           513 => x"a4",
           514 => x"90",
           515 => x"a4",
           516 => x"c8",
           517 => x"a4",
           518 => x"90",
           519 => x"a4",
           520 => x"f3",
           521 => x"a4",
           522 => x"90",
           523 => x"a4",
           524 => x"d6",
           525 => x"a4",
           526 => x"90",
           527 => x"a4",
           528 => x"ab",
           529 => x"a4",
           530 => x"90",
           531 => x"a4",
           532 => x"b5",
           533 => x"a4",
           534 => x"90",
           535 => x"a4",
           536 => x"f7",
           537 => x"a4",
           538 => x"90",
           539 => x"a4",
           540 => x"bd",
           541 => x"a4",
           542 => x"90",
           543 => x"a4",
           544 => x"e3",
           545 => x"a4",
           546 => x"90",
           547 => x"a4",
           548 => x"98",
           549 => x"a4",
           550 => x"90",
           551 => x"a4",
           552 => x"84",
           553 => x"a4",
           554 => x"90",
           555 => x"a4",
           556 => x"f8",
           557 => x"a4",
           558 => x"90",
           559 => x"a4",
           560 => x"e2",
           561 => x"a4",
           562 => x"90",
           563 => x"a4",
           564 => x"c6",
           565 => x"a4",
           566 => x"90",
           567 => x"a4",
           568 => x"ec",
           569 => x"a4",
           570 => x"90",
           571 => x"a4",
           572 => x"90",
           573 => x"a4",
           574 => x"90",
           575 => x"a4",
           576 => x"f3",
           577 => x"a4",
           578 => x"90",
           579 => x"a4",
           580 => x"98",
           581 => x"a4",
           582 => x"90",
           583 => x"a4",
           584 => x"8c",
           585 => x"a4",
           586 => x"90",
           587 => x"a4",
           588 => x"b4",
           589 => x"a4",
           590 => x"90",
           591 => x"a4",
           592 => x"ac",
           593 => x"a4",
           594 => x"90",
           595 => x"a4",
           596 => x"f6",
           597 => x"a4",
           598 => x"90",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"00",
           609 => x"ff",
           610 => x"06",
           611 => x"83",
           612 => x"10",
           613 => x"fc",
           614 => x"51",
           615 => x"80",
           616 => x"ff",
           617 => x"06",
           618 => x"52",
           619 => x"0a",
           620 => x"38",
           621 => x"51",
           622 => x"98",
           623 => x"f4",
           624 => x"80",
           625 => x"05",
           626 => x"0b",
           627 => x"04",
           628 => x"80",
           629 => x"00",
           630 => x"08",
           631 => x"a4",
           632 => x"0d",
           633 => x"08",
           634 => x"82",
           635 => x"fc",
           636 => x"b6",
           637 => x"05",
           638 => x"b6",
           639 => x"05",
           640 => x"cd",
           641 => x"54",
           642 => x"82",
           643 => x"70",
           644 => x"08",
           645 => x"82",
           646 => x"f8",
           647 => x"82",
           648 => x"51",
           649 => x"0d",
           650 => x"0c",
           651 => x"a4",
           652 => x"b6",
           653 => x"3d",
           654 => x"a4",
           655 => x"08",
           656 => x"70",
           657 => x"81",
           658 => x"51",
           659 => x"38",
           660 => x"b6",
           661 => x"05",
           662 => x"38",
           663 => x"0b",
           664 => x"08",
           665 => x"81",
           666 => x"b6",
           667 => x"05",
           668 => x"82",
           669 => x"8c",
           670 => x"0b",
           671 => x"08",
           672 => x"82",
           673 => x"88",
           674 => x"b6",
           675 => x"05",
           676 => x"a4",
           677 => x"08",
           678 => x"f6",
           679 => x"82",
           680 => x"8c",
           681 => x"80",
           682 => x"b6",
           683 => x"05",
           684 => x"90",
           685 => x"98",
           686 => x"b6",
           687 => x"05",
           688 => x"b6",
           689 => x"05",
           690 => x"09",
           691 => x"38",
           692 => x"b6",
           693 => x"05",
           694 => x"39",
           695 => x"08",
           696 => x"82",
           697 => x"f8",
           698 => x"53",
           699 => x"82",
           700 => x"8c",
           701 => x"05",
           702 => x"08",
           703 => x"82",
           704 => x"fc",
           705 => x"05",
           706 => x"08",
           707 => x"ff",
           708 => x"b6",
           709 => x"05",
           710 => x"72",
           711 => x"a4",
           712 => x"08",
           713 => x"a4",
           714 => x"0c",
           715 => x"a4",
           716 => x"08",
           717 => x"0c",
           718 => x"82",
           719 => x"04",
           720 => x"08",
           721 => x"a4",
           722 => x"0d",
           723 => x"b6",
           724 => x"05",
           725 => x"a4",
           726 => x"08",
           727 => x"08",
           728 => x"fe",
           729 => x"b6",
           730 => x"05",
           731 => x"a4",
           732 => x"70",
           733 => x"08",
           734 => x"82",
           735 => x"fc",
           736 => x"82",
           737 => x"8c",
           738 => x"82",
           739 => x"e0",
           740 => x"51",
           741 => x"3f",
           742 => x"08",
           743 => x"a4",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"88",
           748 => x"51",
           749 => x"34",
           750 => x"08",
           751 => x"70",
           752 => x"0c",
           753 => x"0d",
           754 => x"0c",
           755 => x"a4",
           756 => x"b6",
           757 => x"3d",
           758 => x"a4",
           759 => x"70",
           760 => x"08",
           761 => x"82",
           762 => x"fc",
           763 => x"82",
           764 => x"8c",
           765 => x"82",
           766 => x"88",
           767 => x"54",
           768 => x"b6",
           769 => x"82",
           770 => x"f8",
           771 => x"b6",
           772 => x"05",
           773 => x"b6",
           774 => x"54",
           775 => x"82",
           776 => x"04",
           777 => x"08",
           778 => x"a4",
           779 => x"0d",
           780 => x"b6",
           781 => x"05",
           782 => x"a4",
           783 => x"08",
           784 => x"8c",
           785 => x"b6",
           786 => x"05",
           787 => x"33",
           788 => x"70",
           789 => x"81",
           790 => x"51",
           791 => x"80",
           792 => x"ff",
           793 => x"a4",
           794 => x"0c",
           795 => x"82",
           796 => x"8c",
           797 => x"72",
           798 => x"82",
           799 => x"f8",
           800 => x"81",
           801 => x"72",
           802 => x"fa",
           803 => x"a4",
           804 => x"08",
           805 => x"b6",
           806 => x"05",
           807 => x"a4",
           808 => x"22",
           809 => x"51",
           810 => x"2e",
           811 => x"82",
           812 => x"f8",
           813 => x"af",
           814 => x"fc",
           815 => x"a4",
           816 => x"33",
           817 => x"26",
           818 => x"82",
           819 => x"f8",
           820 => x"72",
           821 => x"81",
           822 => x"38",
           823 => x"08",
           824 => x"70",
           825 => x"98",
           826 => x"53",
           827 => x"82",
           828 => x"e4",
           829 => x"83",
           830 => x"32",
           831 => x"51",
           832 => x"72",
           833 => x"38",
           834 => x"08",
           835 => x"70",
           836 => x"51",
           837 => x"b6",
           838 => x"05",
           839 => x"39",
           840 => x"08",
           841 => x"70",
           842 => x"98",
           843 => x"83",
           844 => x"73",
           845 => x"51",
           846 => x"53",
           847 => x"a4",
           848 => x"34",
           849 => x"08",
           850 => x"54",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"82",
           855 => x"e8",
           856 => x"b6",
           857 => x"05",
           858 => x"2b",
           859 => x"51",
           860 => x"80",
           861 => x"80",
           862 => x"b6",
           863 => x"05",
           864 => x"a4",
           865 => x"22",
           866 => x"70",
           867 => x"51",
           868 => x"db",
           869 => x"a4",
           870 => x"33",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"b6",
           876 => x"05",
           877 => x"39",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"9d",
           883 => x"a4",
           884 => x"33",
           885 => x"70",
           886 => x"51",
           887 => x"38",
           888 => x"b6",
           889 => x"05",
           890 => x"a4",
           891 => x"33",
           892 => x"b6",
           893 => x"05",
           894 => x"b6",
           895 => x"05",
           896 => x"26",
           897 => x"82",
           898 => x"c4",
           899 => x"82",
           900 => x"88",
           901 => x"51",
           902 => x"72",
           903 => x"a4",
           904 => x"22",
           905 => x"51",
           906 => x"b6",
           907 => x"05",
           908 => x"a4",
           909 => x"22",
           910 => x"51",
           911 => x"b6",
           912 => x"05",
           913 => x"39",
           914 => x"08",
           915 => x"70",
           916 => x"51",
           917 => x"b6",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"51",
           923 => x"b6",
           924 => x"05",
           925 => x"39",
           926 => x"08",
           927 => x"70",
           928 => x"53",
           929 => x"a4",
           930 => x"23",
           931 => x"b6",
           932 => x"05",
           933 => x"39",
           934 => x"08",
           935 => x"70",
           936 => x"53",
           937 => x"a4",
           938 => x"23",
           939 => x"bf",
           940 => x"a4",
           941 => x"34",
           942 => x"08",
           943 => x"ff",
           944 => x"72",
           945 => x"08",
           946 => x"80",
           947 => x"b6",
           948 => x"05",
           949 => x"39",
           950 => x"08",
           951 => x"82",
           952 => x"90",
           953 => x"05",
           954 => x"08",
           955 => x"70",
           956 => x"72",
           957 => x"08",
           958 => x"82",
           959 => x"ec",
           960 => x"11",
           961 => x"82",
           962 => x"ec",
           963 => x"ef",
           964 => x"a4",
           965 => x"08",
           966 => x"08",
           967 => x"84",
           968 => x"a4",
           969 => x"0c",
           970 => x"b6",
           971 => x"05",
           972 => x"a4",
           973 => x"22",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"82",
           978 => x"e8",
           979 => x"98",
           980 => x"98",
           981 => x"b6",
           982 => x"05",
           983 => x"a2",
           984 => x"b6",
           985 => x"72",
           986 => x"08",
           987 => x"99",
           988 => x"a4",
           989 => x"08",
           990 => x"3f",
           991 => x"08",
           992 => x"b6",
           993 => x"05",
           994 => x"a4",
           995 => x"22",
           996 => x"a4",
           997 => x"22",
           998 => x"54",
           999 => x"b6",
          1000 => x"05",
          1001 => x"39",
          1002 => x"08",
          1003 => x"82",
          1004 => x"90",
          1005 => x"05",
          1006 => x"08",
          1007 => x"70",
          1008 => x"a4",
          1009 => x"0c",
          1010 => x"08",
          1011 => x"70",
          1012 => x"81",
          1013 => x"51",
          1014 => x"2e",
          1015 => x"b6",
          1016 => x"05",
          1017 => x"2b",
          1018 => x"2c",
          1019 => x"a4",
          1020 => x"08",
          1021 => x"c1",
          1022 => x"98",
          1023 => x"82",
          1024 => x"f4",
          1025 => x"39",
          1026 => x"08",
          1027 => x"51",
          1028 => x"82",
          1029 => x"53",
          1030 => x"a4",
          1031 => x"23",
          1032 => x"08",
          1033 => x"53",
          1034 => x"08",
          1035 => x"73",
          1036 => x"54",
          1037 => x"a4",
          1038 => x"23",
          1039 => x"82",
          1040 => x"e4",
          1041 => x"82",
          1042 => x"06",
          1043 => x"72",
          1044 => x"38",
          1045 => x"08",
          1046 => x"82",
          1047 => x"90",
          1048 => x"05",
          1049 => x"08",
          1050 => x"70",
          1051 => x"a4",
          1052 => x"0c",
          1053 => x"82",
          1054 => x"90",
          1055 => x"b6",
          1056 => x"05",
          1057 => x"82",
          1058 => x"90",
          1059 => x"08",
          1060 => x"08",
          1061 => x"53",
          1062 => x"08",
          1063 => x"82",
          1064 => x"fc",
          1065 => x"b6",
          1066 => x"05",
          1067 => x"a4",
          1068 => x"a4",
          1069 => x"22",
          1070 => x"51",
          1071 => x"b6",
          1072 => x"05",
          1073 => x"a4",
          1074 => x"08",
          1075 => x"a4",
          1076 => x"0c",
          1077 => x"08",
          1078 => x"70",
          1079 => x"51",
          1080 => x"b6",
          1081 => x"05",
          1082 => x"39",
          1083 => x"b6",
          1084 => x"05",
          1085 => x"82",
          1086 => x"e4",
          1087 => x"80",
          1088 => x"53",
          1089 => x"a4",
          1090 => x"23",
          1091 => x"82",
          1092 => x"f8",
          1093 => x"0b",
          1094 => x"08",
          1095 => x"82",
          1096 => x"e4",
          1097 => x"82",
          1098 => x"06",
          1099 => x"72",
          1100 => x"38",
          1101 => x"08",
          1102 => x"82",
          1103 => x"90",
          1104 => x"05",
          1105 => x"08",
          1106 => x"70",
          1107 => x"a4",
          1108 => x"0c",
          1109 => x"82",
          1110 => x"90",
          1111 => x"b6",
          1112 => x"05",
          1113 => x"82",
          1114 => x"90",
          1115 => x"08",
          1116 => x"08",
          1117 => x"53",
          1118 => x"08",
          1119 => x"82",
          1120 => x"fc",
          1121 => x"b6",
          1122 => x"05",
          1123 => x"06",
          1124 => x"82",
          1125 => x"e4",
          1126 => x"b6",
          1127 => x"b6",
          1128 => x"05",
          1129 => x"a4",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"55",
          1135 => x"54",
          1136 => x"3f",
          1137 => x"08",
          1138 => x"34",
          1139 => x"08",
          1140 => x"82",
          1141 => x"d4",
          1142 => x"b6",
          1143 => x"05",
          1144 => x"51",
          1145 => x"27",
          1146 => x"b6",
          1147 => x"05",
          1148 => x"33",
          1149 => x"a4",
          1150 => x"33",
          1151 => x"11",
          1152 => x"72",
          1153 => x"08",
          1154 => x"97",
          1155 => x"a4",
          1156 => x"08",
          1157 => x"b0",
          1158 => x"72",
          1159 => x"08",
          1160 => x"82",
          1161 => x"d4",
          1162 => x"82",
          1163 => x"d0",
          1164 => x"34",
          1165 => x"08",
          1166 => x"81",
          1167 => x"a4",
          1168 => x"0c",
          1169 => x"08",
          1170 => x"70",
          1171 => x"a4",
          1172 => x"08",
          1173 => x"ab",
          1174 => x"98",
          1175 => x"b6",
          1176 => x"05",
          1177 => x"b6",
          1178 => x"05",
          1179 => x"84",
          1180 => x"39",
          1181 => x"08",
          1182 => x"82",
          1183 => x"55",
          1184 => x"70",
          1185 => x"53",
          1186 => x"a4",
          1187 => x"34",
          1188 => x"08",
          1189 => x"70",
          1190 => x"53",
          1191 => x"94",
          1192 => x"a4",
          1193 => x"22",
          1194 => x"53",
          1195 => x"a4",
          1196 => x"23",
          1197 => x"08",
          1198 => x"70",
          1199 => x"81",
          1200 => x"53",
          1201 => x"80",
          1202 => x"b6",
          1203 => x"05",
          1204 => x"2b",
          1205 => x"08",
          1206 => x"82",
          1207 => x"cc",
          1208 => x"2c",
          1209 => x"08",
          1210 => x"82",
          1211 => x"f4",
          1212 => x"53",
          1213 => x"09",
          1214 => x"38",
          1215 => x"08",
          1216 => x"fe",
          1217 => x"82",
          1218 => x"c8",
          1219 => x"39",
          1220 => x"08",
          1221 => x"ff",
          1222 => x"82",
          1223 => x"c8",
          1224 => x"b6",
          1225 => x"05",
          1226 => x"a4",
          1227 => x"23",
          1228 => x"08",
          1229 => x"70",
          1230 => x"81",
          1231 => x"53",
          1232 => x"80",
          1233 => x"b6",
          1234 => x"05",
          1235 => x"2b",
          1236 => x"82",
          1237 => x"fc",
          1238 => x"51",
          1239 => x"74",
          1240 => x"82",
          1241 => x"e4",
          1242 => x"f7",
          1243 => x"72",
          1244 => x"08",
          1245 => x"9d",
          1246 => x"a4",
          1247 => x"33",
          1248 => x"a4",
          1249 => x"33",
          1250 => x"54",
          1251 => x"b6",
          1252 => x"05",
          1253 => x"a4",
          1254 => x"22",
          1255 => x"70",
          1256 => x"51",
          1257 => x"2e",
          1258 => x"b6",
          1259 => x"05",
          1260 => x"2b",
          1261 => x"70",
          1262 => x"88",
          1263 => x"51",
          1264 => x"54",
          1265 => x"08",
          1266 => x"70",
          1267 => x"53",
          1268 => x"a4",
          1269 => x"23",
          1270 => x"b6",
          1271 => x"05",
          1272 => x"2b",
          1273 => x"70",
          1274 => x"88",
          1275 => x"51",
          1276 => x"54",
          1277 => x"08",
          1278 => x"70",
          1279 => x"53",
          1280 => x"a4",
          1281 => x"23",
          1282 => x"08",
          1283 => x"70",
          1284 => x"51",
          1285 => x"38",
          1286 => x"08",
          1287 => x"ff",
          1288 => x"72",
          1289 => x"08",
          1290 => x"73",
          1291 => x"90",
          1292 => x"80",
          1293 => x"38",
          1294 => x"08",
          1295 => x"52",
          1296 => x"ee",
          1297 => x"82",
          1298 => x"e4",
          1299 => x"81",
          1300 => x"06",
          1301 => x"72",
          1302 => x"38",
          1303 => x"08",
          1304 => x"52",
          1305 => x"ca",
          1306 => x"39",
          1307 => x"08",
          1308 => x"70",
          1309 => x"81",
          1310 => x"53",
          1311 => x"90",
          1312 => x"a4",
          1313 => x"08",
          1314 => x"8a",
          1315 => x"39",
          1316 => x"08",
          1317 => x"70",
          1318 => x"81",
          1319 => x"53",
          1320 => x"8e",
          1321 => x"a4",
          1322 => x"08",
          1323 => x"8a",
          1324 => x"b6",
          1325 => x"05",
          1326 => x"2a",
          1327 => x"51",
          1328 => x"80",
          1329 => x"82",
          1330 => x"88",
          1331 => x"b0",
          1332 => x"3f",
          1333 => x"08",
          1334 => x"53",
          1335 => x"09",
          1336 => x"38",
          1337 => x"08",
          1338 => x"52",
          1339 => x"08",
          1340 => x"51",
          1341 => x"82",
          1342 => x"e4",
          1343 => x"88",
          1344 => x"06",
          1345 => x"72",
          1346 => x"38",
          1347 => x"08",
          1348 => x"ff",
          1349 => x"72",
          1350 => x"08",
          1351 => x"73",
          1352 => x"90",
          1353 => x"80",
          1354 => x"38",
          1355 => x"08",
          1356 => x"52",
          1357 => x"fa",
          1358 => x"82",
          1359 => x"e4",
          1360 => x"83",
          1361 => x"06",
          1362 => x"72",
          1363 => x"38",
          1364 => x"08",
          1365 => x"ff",
          1366 => x"72",
          1367 => x"08",
          1368 => x"73",
          1369 => x"98",
          1370 => x"80",
          1371 => x"38",
          1372 => x"08",
          1373 => x"52",
          1374 => x"b6",
          1375 => x"82",
          1376 => x"e4",
          1377 => x"87",
          1378 => x"06",
          1379 => x"72",
          1380 => x"b6",
          1381 => x"05",
          1382 => x"54",
          1383 => x"b6",
          1384 => x"05",
          1385 => x"2b",
          1386 => x"51",
          1387 => x"25",
          1388 => x"b6",
          1389 => x"05",
          1390 => x"51",
          1391 => x"d2",
          1392 => x"a4",
          1393 => x"33",
          1394 => x"e3",
          1395 => x"06",
          1396 => x"b6",
          1397 => x"05",
          1398 => x"b6",
          1399 => x"05",
          1400 => x"ce",
          1401 => x"39",
          1402 => x"08",
          1403 => x"53",
          1404 => x"2e",
          1405 => x"80",
          1406 => x"b6",
          1407 => x"05",
          1408 => x"51",
          1409 => x"b6",
          1410 => x"05",
          1411 => x"ff",
          1412 => x"72",
          1413 => x"2e",
          1414 => x"82",
          1415 => x"88",
          1416 => x"82",
          1417 => x"fc",
          1418 => x"33",
          1419 => x"a4",
          1420 => x"08",
          1421 => x"b6",
          1422 => x"05",
          1423 => x"f2",
          1424 => x"39",
          1425 => x"08",
          1426 => x"53",
          1427 => x"2e",
          1428 => x"80",
          1429 => x"b6",
          1430 => x"05",
          1431 => x"51",
          1432 => x"b6",
          1433 => x"05",
          1434 => x"ff",
          1435 => x"72",
          1436 => x"2e",
          1437 => x"82",
          1438 => x"88",
          1439 => x"82",
          1440 => x"fc",
          1441 => x"33",
          1442 => x"a6",
          1443 => x"a4",
          1444 => x"08",
          1445 => x"b6",
          1446 => x"05",
          1447 => x"39",
          1448 => x"08",
          1449 => x"82",
          1450 => x"a9",
          1451 => x"a4",
          1452 => x"08",
          1453 => x"a4",
          1454 => x"08",
          1455 => x"b6",
          1456 => x"05",
          1457 => x"a4",
          1458 => x"08",
          1459 => x"53",
          1460 => x"cc",
          1461 => x"a4",
          1462 => x"22",
          1463 => x"70",
          1464 => x"51",
          1465 => x"2e",
          1466 => x"82",
          1467 => x"ec",
          1468 => x"11",
          1469 => x"82",
          1470 => x"ec",
          1471 => x"90",
          1472 => x"2c",
          1473 => x"73",
          1474 => x"82",
          1475 => x"88",
          1476 => x"a0",
          1477 => x"3f",
          1478 => x"b6",
          1479 => x"05",
          1480 => x"b6",
          1481 => x"05",
          1482 => x"86",
          1483 => x"82",
          1484 => x"e4",
          1485 => x"b7",
          1486 => x"a4",
          1487 => x"33",
          1488 => x"2e",
          1489 => x"a8",
          1490 => x"82",
          1491 => x"e4",
          1492 => x"0b",
          1493 => x"08",
          1494 => x"80",
          1495 => x"a4",
          1496 => x"34",
          1497 => x"b6",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"52",
          1502 => x"08",
          1503 => x"51",
          1504 => x"e9",
          1505 => x"b6",
          1506 => x"05",
          1507 => x"08",
          1508 => x"a4",
          1509 => x"0c",
          1510 => x"b6",
          1511 => x"05",
          1512 => x"98",
          1513 => x"0d",
          1514 => x"0c",
          1515 => x"a4",
          1516 => x"b6",
          1517 => x"3d",
          1518 => x"e8",
          1519 => x"b6",
          1520 => x"05",
          1521 => x"b6",
          1522 => x"05",
          1523 => x"dd",
          1524 => x"98",
          1525 => x"b6",
          1526 => x"85",
          1527 => x"b6",
          1528 => x"82",
          1529 => x"02",
          1530 => x"0c",
          1531 => x"80",
          1532 => x"a4",
          1533 => x"0c",
          1534 => x"08",
          1535 => x"70",
          1536 => x"81",
          1537 => x"06",
          1538 => x"51",
          1539 => x"2e",
          1540 => x"0b",
          1541 => x"08",
          1542 => x"81",
          1543 => x"b6",
          1544 => x"05",
          1545 => x"33",
          1546 => x"08",
          1547 => x"81",
          1548 => x"a4",
          1549 => x"0c",
          1550 => x"b6",
          1551 => x"05",
          1552 => x"ff",
          1553 => x"80",
          1554 => x"82",
          1555 => x"82",
          1556 => x"53",
          1557 => x"08",
          1558 => x"52",
          1559 => x"51",
          1560 => x"82",
          1561 => x"53",
          1562 => x"ff",
          1563 => x"0b",
          1564 => x"08",
          1565 => x"ff",
          1566 => x"cd",
          1567 => x"cd",
          1568 => x"53",
          1569 => x"13",
          1570 => x"2d",
          1571 => x"08",
          1572 => x"2e",
          1573 => x"0b",
          1574 => x"08",
          1575 => x"82",
          1576 => x"f8",
          1577 => x"82",
          1578 => x"f4",
          1579 => x"82",
          1580 => x"f4",
          1581 => x"b6",
          1582 => x"3d",
          1583 => x"a4",
          1584 => x"b6",
          1585 => x"82",
          1586 => x"fb",
          1587 => x"0b",
          1588 => x"08",
          1589 => x"82",
          1590 => x"8c",
          1591 => x"11",
          1592 => x"2a",
          1593 => x"70",
          1594 => x"51",
          1595 => x"72",
          1596 => x"38",
          1597 => x"b6",
          1598 => x"05",
          1599 => x"39",
          1600 => x"08",
          1601 => x"53",
          1602 => x"b6",
          1603 => x"05",
          1604 => x"82",
          1605 => x"88",
          1606 => x"72",
          1607 => x"08",
          1608 => x"72",
          1609 => x"53",
          1610 => x"b6",
          1611 => x"a4",
          1612 => x"08",
          1613 => x"08",
          1614 => x"53",
          1615 => x"08",
          1616 => x"52",
          1617 => x"51",
          1618 => x"82",
          1619 => x"53",
          1620 => x"ff",
          1621 => x"0b",
          1622 => x"08",
          1623 => x"ff",
          1624 => x"b6",
          1625 => x"05",
          1626 => x"b6",
          1627 => x"05",
          1628 => x"b6",
          1629 => x"05",
          1630 => x"98",
          1631 => x"0d",
          1632 => x"0c",
          1633 => x"a4",
          1634 => x"b6",
          1635 => x"3d",
          1636 => x"ec",
          1637 => x"b6",
          1638 => x"05",
          1639 => x"3f",
          1640 => x"08",
          1641 => x"98",
          1642 => x"3d",
          1643 => x"a4",
          1644 => x"b6",
          1645 => x"82",
          1646 => x"fb",
          1647 => x"b6",
          1648 => x"05",
          1649 => x"33",
          1650 => x"70",
          1651 => x"81",
          1652 => x"51",
          1653 => x"80",
          1654 => x"ff",
          1655 => x"a4",
          1656 => x"0c",
          1657 => x"82",
          1658 => x"8c",
          1659 => x"11",
          1660 => x"2a",
          1661 => x"51",
          1662 => x"72",
          1663 => x"db",
          1664 => x"a4",
          1665 => x"08",
          1666 => x"08",
          1667 => x"54",
          1668 => x"08",
          1669 => x"25",
          1670 => x"b6",
          1671 => x"05",
          1672 => x"70",
          1673 => x"08",
          1674 => x"52",
          1675 => x"72",
          1676 => x"08",
          1677 => x"0c",
          1678 => x"08",
          1679 => x"8c",
          1680 => x"05",
          1681 => x"82",
          1682 => x"88",
          1683 => x"82",
          1684 => x"fc",
          1685 => x"53",
          1686 => x"82",
          1687 => x"8c",
          1688 => x"b6",
          1689 => x"05",
          1690 => x"b6",
          1691 => x"05",
          1692 => x"ff",
          1693 => x"12",
          1694 => x"54",
          1695 => x"b6",
          1696 => x"72",
          1697 => x"b6",
          1698 => x"05",
          1699 => x"08",
          1700 => x"12",
          1701 => x"a4",
          1702 => x"08",
          1703 => x"a4",
          1704 => x"0c",
          1705 => x"39",
          1706 => x"b6",
          1707 => x"05",
          1708 => x"a4",
          1709 => x"08",
          1710 => x"0c",
          1711 => x"82",
          1712 => x"04",
          1713 => x"08",
          1714 => x"a4",
          1715 => x"0d",
          1716 => x"08",
          1717 => x"85",
          1718 => x"81",
          1719 => x"06",
          1720 => x"52",
          1721 => x"8d",
          1722 => x"82",
          1723 => x"f8",
          1724 => x"94",
          1725 => x"a4",
          1726 => x"08",
          1727 => x"70",
          1728 => x"81",
          1729 => x"51",
          1730 => x"2e",
          1731 => x"82",
          1732 => x"88",
          1733 => x"b6",
          1734 => x"05",
          1735 => x"85",
          1736 => x"ff",
          1737 => x"52",
          1738 => x"34",
          1739 => x"08",
          1740 => x"8c",
          1741 => x"05",
          1742 => x"82",
          1743 => x"88",
          1744 => x"11",
          1745 => x"b6",
          1746 => x"05",
          1747 => x"52",
          1748 => x"82",
          1749 => x"88",
          1750 => x"11",
          1751 => x"2a",
          1752 => x"51",
          1753 => x"71",
          1754 => x"d7",
          1755 => x"a4",
          1756 => x"08",
          1757 => x"33",
          1758 => x"08",
          1759 => x"51",
          1760 => x"a4",
          1761 => x"08",
          1762 => x"b6",
          1763 => x"05",
          1764 => x"a4",
          1765 => x"08",
          1766 => x"12",
          1767 => x"07",
          1768 => x"85",
          1769 => x"0b",
          1770 => x"08",
          1771 => x"81",
          1772 => x"b6",
          1773 => x"05",
          1774 => x"81",
          1775 => x"52",
          1776 => x"82",
          1777 => x"88",
          1778 => x"b6",
          1779 => x"05",
          1780 => x"11",
          1781 => x"71",
          1782 => x"98",
          1783 => x"b6",
          1784 => x"05",
          1785 => x"b6",
          1786 => x"05",
          1787 => x"80",
          1788 => x"b6",
          1789 => x"05",
          1790 => x"a4",
          1791 => x"0c",
          1792 => x"08",
          1793 => x"85",
          1794 => x"b6",
          1795 => x"05",
          1796 => x"b6",
          1797 => x"05",
          1798 => x"09",
          1799 => x"38",
          1800 => x"08",
          1801 => x"90",
          1802 => x"82",
          1803 => x"ec",
          1804 => x"39",
          1805 => x"08",
          1806 => x"a0",
          1807 => x"82",
          1808 => x"ec",
          1809 => x"b6",
          1810 => x"05",
          1811 => x"b6",
          1812 => x"05",
          1813 => x"34",
          1814 => x"b6",
          1815 => x"05",
          1816 => x"82",
          1817 => x"88",
          1818 => x"11",
          1819 => x"8c",
          1820 => x"b6",
          1821 => x"05",
          1822 => x"ff",
          1823 => x"b6",
          1824 => x"05",
          1825 => x"52",
          1826 => x"08",
          1827 => x"82",
          1828 => x"89",
          1829 => x"b6",
          1830 => x"82",
          1831 => x"02",
          1832 => x"0c",
          1833 => x"82",
          1834 => x"88",
          1835 => x"b6",
          1836 => x"05",
          1837 => x"a4",
          1838 => x"08",
          1839 => x"08",
          1840 => x"82",
          1841 => x"90",
          1842 => x"2e",
          1843 => x"82",
          1844 => x"f8",
          1845 => x"b6",
          1846 => x"05",
          1847 => x"ac",
          1848 => x"a4",
          1849 => x"08",
          1850 => x"08",
          1851 => x"05",
          1852 => x"a4",
          1853 => x"08",
          1854 => x"90",
          1855 => x"a4",
          1856 => x"08",
          1857 => x"08",
          1858 => x"05",
          1859 => x"08",
          1860 => x"82",
          1861 => x"f8",
          1862 => x"b6",
          1863 => x"05",
          1864 => x"b6",
          1865 => x"05",
          1866 => x"a4",
          1867 => x"08",
          1868 => x"b6",
          1869 => x"05",
          1870 => x"a4",
          1871 => x"08",
          1872 => x"b6",
          1873 => x"05",
          1874 => x"a4",
          1875 => x"08",
          1876 => x"9c",
          1877 => x"a4",
          1878 => x"08",
          1879 => x"b6",
          1880 => x"05",
          1881 => x"a4",
          1882 => x"08",
          1883 => x"b6",
          1884 => x"05",
          1885 => x"a4",
          1886 => x"08",
          1887 => x"08",
          1888 => x"53",
          1889 => x"71",
          1890 => x"39",
          1891 => x"08",
          1892 => x"81",
          1893 => x"a4",
          1894 => x"0c",
          1895 => x"08",
          1896 => x"ff",
          1897 => x"a4",
          1898 => x"0c",
          1899 => x"08",
          1900 => x"80",
          1901 => x"82",
          1902 => x"f8",
          1903 => x"70",
          1904 => x"a4",
          1905 => x"08",
          1906 => x"b6",
          1907 => x"05",
          1908 => x"a4",
          1909 => x"08",
          1910 => x"71",
          1911 => x"a4",
          1912 => x"08",
          1913 => x"b6",
          1914 => x"05",
          1915 => x"39",
          1916 => x"08",
          1917 => x"70",
          1918 => x"0c",
          1919 => x"0d",
          1920 => x"0c",
          1921 => x"a4",
          1922 => x"b6",
          1923 => x"3d",
          1924 => x"a4",
          1925 => x"08",
          1926 => x"08",
          1927 => x"82",
          1928 => x"fc",
          1929 => x"71",
          1930 => x"a4",
          1931 => x"08",
          1932 => x"b6",
          1933 => x"05",
          1934 => x"ff",
          1935 => x"70",
          1936 => x"38",
          1937 => x"b6",
          1938 => x"05",
          1939 => x"82",
          1940 => x"fc",
          1941 => x"b6",
          1942 => x"05",
          1943 => x"a4",
          1944 => x"08",
          1945 => x"b6",
          1946 => x"84",
          1947 => x"b6",
          1948 => x"82",
          1949 => x"02",
          1950 => x"0c",
          1951 => x"82",
          1952 => x"88",
          1953 => x"b6",
          1954 => x"05",
          1955 => x"a4",
          1956 => x"08",
          1957 => x"82",
          1958 => x"8c",
          1959 => x"05",
          1960 => x"08",
          1961 => x"82",
          1962 => x"fc",
          1963 => x"51",
          1964 => x"82",
          1965 => x"fc",
          1966 => x"05",
          1967 => x"08",
          1968 => x"70",
          1969 => x"51",
          1970 => x"84",
          1971 => x"39",
          1972 => x"08",
          1973 => x"70",
          1974 => x"0c",
          1975 => x"0d",
          1976 => x"0c",
          1977 => x"a4",
          1978 => x"b6",
          1979 => x"3d",
          1980 => x"a4",
          1981 => x"08",
          1982 => x"08",
          1983 => x"82",
          1984 => x"8c",
          1985 => x"b6",
          1986 => x"05",
          1987 => x"a4",
          1988 => x"08",
          1989 => x"e5",
          1990 => x"a4",
          1991 => x"08",
          1992 => x"b6",
          1993 => x"05",
          1994 => x"a4",
          1995 => x"08",
          1996 => x"b6",
          1997 => x"05",
          1998 => x"a4",
          1999 => x"08",
          2000 => x"38",
          2001 => x"08",
          2002 => x"51",
          2003 => x"b6",
          2004 => x"05",
          2005 => x"82",
          2006 => x"f8",
          2007 => x"b6",
          2008 => x"05",
          2009 => x"71",
          2010 => x"b6",
          2011 => x"05",
          2012 => x"82",
          2013 => x"fc",
          2014 => x"ad",
          2015 => x"a4",
          2016 => x"08",
          2017 => x"98",
          2018 => x"3d",
          2019 => x"a4",
          2020 => x"b6",
          2021 => x"82",
          2022 => x"fd",
          2023 => x"b6",
          2024 => x"05",
          2025 => x"81",
          2026 => x"b6",
          2027 => x"05",
          2028 => x"33",
          2029 => x"08",
          2030 => x"81",
          2031 => x"a4",
          2032 => x"0c",
          2033 => x"08",
          2034 => x"70",
          2035 => x"ff",
          2036 => x"54",
          2037 => x"2e",
          2038 => x"ce",
          2039 => x"a4",
          2040 => x"08",
          2041 => x"82",
          2042 => x"88",
          2043 => x"05",
          2044 => x"08",
          2045 => x"70",
          2046 => x"51",
          2047 => x"38",
          2048 => x"b6",
          2049 => x"05",
          2050 => x"39",
          2051 => x"08",
          2052 => x"ff",
          2053 => x"a4",
          2054 => x"0c",
          2055 => x"08",
          2056 => x"80",
          2057 => x"ff",
          2058 => x"b6",
          2059 => x"05",
          2060 => x"80",
          2061 => x"b6",
          2062 => x"05",
          2063 => x"52",
          2064 => x"38",
          2065 => x"b6",
          2066 => x"05",
          2067 => x"39",
          2068 => x"08",
          2069 => x"ff",
          2070 => x"a4",
          2071 => x"0c",
          2072 => x"08",
          2073 => x"70",
          2074 => x"70",
          2075 => x"0b",
          2076 => x"08",
          2077 => x"ae",
          2078 => x"a4",
          2079 => x"08",
          2080 => x"b6",
          2081 => x"05",
          2082 => x"72",
          2083 => x"82",
          2084 => x"fc",
          2085 => x"55",
          2086 => x"8a",
          2087 => x"82",
          2088 => x"fc",
          2089 => x"b6",
          2090 => x"05",
          2091 => x"98",
          2092 => x"0d",
          2093 => x"0c",
          2094 => x"a4",
          2095 => x"b6",
          2096 => x"3d",
          2097 => x"a4",
          2098 => x"08",
          2099 => x"08",
          2100 => x"82",
          2101 => x"8c",
          2102 => x"38",
          2103 => x"b6",
          2104 => x"05",
          2105 => x"39",
          2106 => x"08",
          2107 => x"52",
          2108 => x"b6",
          2109 => x"05",
          2110 => x"82",
          2111 => x"f8",
          2112 => x"81",
          2113 => x"51",
          2114 => x"9f",
          2115 => x"a4",
          2116 => x"08",
          2117 => x"b6",
          2118 => x"05",
          2119 => x"a4",
          2120 => x"08",
          2121 => x"38",
          2122 => x"82",
          2123 => x"f8",
          2124 => x"05",
          2125 => x"08",
          2126 => x"82",
          2127 => x"f8",
          2128 => x"b6",
          2129 => x"05",
          2130 => x"82",
          2131 => x"fc",
          2132 => x"82",
          2133 => x"fc",
          2134 => x"b6",
          2135 => x"3d",
          2136 => x"a4",
          2137 => x"b6",
          2138 => x"82",
          2139 => x"fe",
          2140 => x"b6",
          2141 => x"05",
          2142 => x"a4",
          2143 => x"0c",
          2144 => x"08",
          2145 => x"80",
          2146 => x"38",
          2147 => x"08",
          2148 => x"81",
          2149 => x"a4",
          2150 => x"0c",
          2151 => x"08",
          2152 => x"ff",
          2153 => x"a4",
          2154 => x"0c",
          2155 => x"08",
          2156 => x"80",
          2157 => x"82",
          2158 => x"8c",
          2159 => x"70",
          2160 => x"08",
          2161 => x"52",
          2162 => x"34",
          2163 => x"08",
          2164 => x"81",
          2165 => x"a4",
          2166 => x"0c",
          2167 => x"82",
          2168 => x"88",
          2169 => x"82",
          2170 => x"51",
          2171 => x"82",
          2172 => x"04",
          2173 => x"08",
          2174 => x"a4",
          2175 => x"0d",
          2176 => x"b6",
          2177 => x"05",
          2178 => x"a4",
          2179 => x"08",
          2180 => x"38",
          2181 => x"08",
          2182 => x"30",
          2183 => x"08",
          2184 => x"80",
          2185 => x"a4",
          2186 => x"0c",
          2187 => x"08",
          2188 => x"8a",
          2189 => x"82",
          2190 => x"f4",
          2191 => x"b6",
          2192 => x"05",
          2193 => x"a4",
          2194 => x"0c",
          2195 => x"08",
          2196 => x"80",
          2197 => x"82",
          2198 => x"8c",
          2199 => x"82",
          2200 => x"8c",
          2201 => x"0b",
          2202 => x"08",
          2203 => x"82",
          2204 => x"fc",
          2205 => x"38",
          2206 => x"b6",
          2207 => x"05",
          2208 => x"a4",
          2209 => x"08",
          2210 => x"08",
          2211 => x"80",
          2212 => x"a4",
          2213 => x"08",
          2214 => x"a4",
          2215 => x"08",
          2216 => x"3f",
          2217 => x"08",
          2218 => x"a4",
          2219 => x"0c",
          2220 => x"a4",
          2221 => x"08",
          2222 => x"38",
          2223 => x"08",
          2224 => x"30",
          2225 => x"08",
          2226 => x"82",
          2227 => x"f8",
          2228 => x"82",
          2229 => x"54",
          2230 => x"82",
          2231 => x"04",
          2232 => x"08",
          2233 => x"a4",
          2234 => x"0d",
          2235 => x"b6",
          2236 => x"05",
          2237 => x"a4",
          2238 => x"08",
          2239 => x"38",
          2240 => x"08",
          2241 => x"30",
          2242 => x"08",
          2243 => x"81",
          2244 => x"a4",
          2245 => x"0c",
          2246 => x"08",
          2247 => x"80",
          2248 => x"82",
          2249 => x"8c",
          2250 => x"82",
          2251 => x"8c",
          2252 => x"53",
          2253 => x"08",
          2254 => x"52",
          2255 => x"08",
          2256 => x"51",
          2257 => x"82",
          2258 => x"70",
          2259 => x"08",
          2260 => x"54",
          2261 => x"08",
          2262 => x"80",
          2263 => x"82",
          2264 => x"f8",
          2265 => x"82",
          2266 => x"f8",
          2267 => x"b6",
          2268 => x"05",
          2269 => x"b6",
          2270 => x"87",
          2271 => x"b6",
          2272 => x"82",
          2273 => x"02",
          2274 => x"0c",
          2275 => x"80",
          2276 => x"a4",
          2277 => x"08",
          2278 => x"a4",
          2279 => x"08",
          2280 => x"3f",
          2281 => x"08",
          2282 => x"98",
          2283 => x"3d",
          2284 => x"a4",
          2285 => x"b6",
          2286 => x"82",
          2287 => x"fd",
          2288 => x"53",
          2289 => x"08",
          2290 => x"52",
          2291 => x"08",
          2292 => x"51",
          2293 => x"b6",
          2294 => x"82",
          2295 => x"54",
          2296 => x"82",
          2297 => x"04",
          2298 => x"08",
          2299 => x"a4",
          2300 => x"0d",
          2301 => x"b6",
          2302 => x"05",
          2303 => x"82",
          2304 => x"f8",
          2305 => x"b6",
          2306 => x"05",
          2307 => x"a4",
          2308 => x"08",
          2309 => x"82",
          2310 => x"fc",
          2311 => x"2e",
          2312 => x"0b",
          2313 => x"08",
          2314 => x"24",
          2315 => x"b6",
          2316 => x"05",
          2317 => x"b6",
          2318 => x"05",
          2319 => x"a4",
          2320 => x"08",
          2321 => x"a4",
          2322 => x"0c",
          2323 => x"82",
          2324 => x"fc",
          2325 => x"2e",
          2326 => x"82",
          2327 => x"8c",
          2328 => x"b6",
          2329 => x"05",
          2330 => x"38",
          2331 => x"08",
          2332 => x"82",
          2333 => x"8c",
          2334 => x"82",
          2335 => x"88",
          2336 => x"b6",
          2337 => x"05",
          2338 => x"a4",
          2339 => x"08",
          2340 => x"a4",
          2341 => x"0c",
          2342 => x"08",
          2343 => x"81",
          2344 => x"a4",
          2345 => x"0c",
          2346 => x"08",
          2347 => x"81",
          2348 => x"a4",
          2349 => x"0c",
          2350 => x"82",
          2351 => x"90",
          2352 => x"2e",
          2353 => x"b6",
          2354 => x"05",
          2355 => x"b6",
          2356 => x"05",
          2357 => x"39",
          2358 => x"08",
          2359 => x"70",
          2360 => x"08",
          2361 => x"51",
          2362 => x"08",
          2363 => x"82",
          2364 => x"85",
          2365 => x"b6",
          2366 => x"82",
          2367 => x"02",
          2368 => x"0c",
          2369 => x"80",
          2370 => x"a4",
          2371 => x"34",
          2372 => x"08",
          2373 => x"53",
          2374 => x"82",
          2375 => x"88",
          2376 => x"08",
          2377 => x"33",
          2378 => x"b6",
          2379 => x"05",
          2380 => x"ff",
          2381 => x"a0",
          2382 => x"06",
          2383 => x"b6",
          2384 => x"05",
          2385 => x"81",
          2386 => x"53",
          2387 => x"b6",
          2388 => x"05",
          2389 => x"ad",
          2390 => x"06",
          2391 => x"0b",
          2392 => x"08",
          2393 => x"82",
          2394 => x"88",
          2395 => x"08",
          2396 => x"0c",
          2397 => x"53",
          2398 => x"b6",
          2399 => x"05",
          2400 => x"a4",
          2401 => x"33",
          2402 => x"2e",
          2403 => x"81",
          2404 => x"b6",
          2405 => x"05",
          2406 => x"81",
          2407 => x"70",
          2408 => x"72",
          2409 => x"a4",
          2410 => x"34",
          2411 => x"08",
          2412 => x"82",
          2413 => x"e8",
          2414 => x"b6",
          2415 => x"05",
          2416 => x"2e",
          2417 => x"b6",
          2418 => x"05",
          2419 => x"2e",
          2420 => x"cd",
          2421 => x"82",
          2422 => x"f4",
          2423 => x"b6",
          2424 => x"05",
          2425 => x"81",
          2426 => x"70",
          2427 => x"72",
          2428 => x"a4",
          2429 => x"34",
          2430 => x"82",
          2431 => x"a4",
          2432 => x"34",
          2433 => x"08",
          2434 => x"70",
          2435 => x"71",
          2436 => x"51",
          2437 => x"82",
          2438 => x"f8",
          2439 => x"fe",
          2440 => x"a4",
          2441 => x"33",
          2442 => x"26",
          2443 => x"0b",
          2444 => x"08",
          2445 => x"83",
          2446 => x"b6",
          2447 => x"05",
          2448 => x"73",
          2449 => x"82",
          2450 => x"f8",
          2451 => x"72",
          2452 => x"38",
          2453 => x"0b",
          2454 => x"08",
          2455 => x"82",
          2456 => x"0b",
          2457 => x"08",
          2458 => x"b2",
          2459 => x"a4",
          2460 => x"33",
          2461 => x"27",
          2462 => x"b6",
          2463 => x"05",
          2464 => x"b9",
          2465 => x"8d",
          2466 => x"82",
          2467 => x"ec",
          2468 => x"a5",
          2469 => x"82",
          2470 => x"f4",
          2471 => x"0b",
          2472 => x"08",
          2473 => x"82",
          2474 => x"f8",
          2475 => x"a0",
          2476 => x"cf",
          2477 => x"a4",
          2478 => x"33",
          2479 => x"73",
          2480 => x"82",
          2481 => x"f8",
          2482 => x"11",
          2483 => x"82",
          2484 => x"f8",
          2485 => x"b6",
          2486 => x"05",
          2487 => x"51",
          2488 => x"b6",
          2489 => x"05",
          2490 => x"a4",
          2491 => x"33",
          2492 => x"27",
          2493 => x"b6",
          2494 => x"05",
          2495 => x"51",
          2496 => x"b6",
          2497 => x"05",
          2498 => x"a4",
          2499 => x"33",
          2500 => x"26",
          2501 => x"0b",
          2502 => x"08",
          2503 => x"81",
          2504 => x"b6",
          2505 => x"05",
          2506 => x"a4",
          2507 => x"33",
          2508 => x"74",
          2509 => x"80",
          2510 => x"a4",
          2511 => x"0c",
          2512 => x"82",
          2513 => x"f4",
          2514 => x"82",
          2515 => x"fc",
          2516 => x"82",
          2517 => x"f8",
          2518 => x"12",
          2519 => x"08",
          2520 => x"82",
          2521 => x"88",
          2522 => x"08",
          2523 => x"0c",
          2524 => x"51",
          2525 => x"72",
          2526 => x"a4",
          2527 => x"34",
          2528 => x"82",
          2529 => x"f0",
          2530 => x"72",
          2531 => x"38",
          2532 => x"08",
          2533 => x"30",
          2534 => x"08",
          2535 => x"82",
          2536 => x"8c",
          2537 => x"b6",
          2538 => x"05",
          2539 => x"53",
          2540 => x"b6",
          2541 => x"05",
          2542 => x"a4",
          2543 => x"08",
          2544 => x"0c",
          2545 => x"82",
          2546 => x"04",
          2547 => x"08",
          2548 => x"a4",
          2549 => x"0d",
          2550 => x"b6",
          2551 => x"05",
          2552 => x"a4",
          2553 => x"08",
          2554 => x"0c",
          2555 => x"08",
          2556 => x"70",
          2557 => x"72",
          2558 => x"82",
          2559 => x"f8",
          2560 => x"81",
          2561 => x"72",
          2562 => x"81",
          2563 => x"82",
          2564 => x"88",
          2565 => x"08",
          2566 => x"0c",
          2567 => x"82",
          2568 => x"f8",
          2569 => x"72",
          2570 => x"81",
          2571 => x"81",
          2572 => x"a4",
          2573 => x"34",
          2574 => x"08",
          2575 => x"70",
          2576 => x"71",
          2577 => x"51",
          2578 => x"82",
          2579 => x"f8",
          2580 => x"b6",
          2581 => x"05",
          2582 => x"b0",
          2583 => x"06",
          2584 => x"82",
          2585 => x"88",
          2586 => x"08",
          2587 => x"0c",
          2588 => x"53",
          2589 => x"b6",
          2590 => x"05",
          2591 => x"a4",
          2592 => x"33",
          2593 => x"08",
          2594 => x"82",
          2595 => x"e8",
          2596 => x"e2",
          2597 => x"82",
          2598 => x"e8",
          2599 => x"f8",
          2600 => x"80",
          2601 => x"0b",
          2602 => x"08",
          2603 => x"82",
          2604 => x"88",
          2605 => x"08",
          2606 => x"0c",
          2607 => x"53",
          2608 => x"b6",
          2609 => x"05",
          2610 => x"39",
          2611 => x"b6",
          2612 => x"05",
          2613 => x"a4",
          2614 => x"08",
          2615 => x"05",
          2616 => x"08",
          2617 => x"33",
          2618 => x"08",
          2619 => x"80",
          2620 => x"b6",
          2621 => x"05",
          2622 => x"a0",
          2623 => x"81",
          2624 => x"a4",
          2625 => x"0c",
          2626 => x"82",
          2627 => x"f8",
          2628 => x"af",
          2629 => x"38",
          2630 => x"08",
          2631 => x"53",
          2632 => x"83",
          2633 => x"80",
          2634 => x"a4",
          2635 => x"0c",
          2636 => x"88",
          2637 => x"a4",
          2638 => x"34",
          2639 => x"b6",
          2640 => x"05",
          2641 => x"73",
          2642 => x"82",
          2643 => x"f8",
          2644 => x"72",
          2645 => x"38",
          2646 => x"0b",
          2647 => x"08",
          2648 => x"82",
          2649 => x"0b",
          2650 => x"08",
          2651 => x"80",
          2652 => x"a4",
          2653 => x"0c",
          2654 => x"08",
          2655 => x"53",
          2656 => x"81",
          2657 => x"b6",
          2658 => x"05",
          2659 => x"e0",
          2660 => x"38",
          2661 => x"08",
          2662 => x"e0",
          2663 => x"72",
          2664 => x"08",
          2665 => x"82",
          2666 => x"f8",
          2667 => x"11",
          2668 => x"82",
          2669 => x"f8",
          2670 => x"b6",
          2671 => x"05",
          2672 => x"73",
          2673 => x"82",
          2674 => x"f8",
          2675 => x"11",
          2676 => x"82",
          2677 => x"f8",
          2678 => x"b6",
          2679 => x"05",
          2680 => x"89",
          2681 => x"80",
          2682 => x"a4",
          2683 => x"0c",
          2684 => x"82",
          2685 => x"f8",
          2686 => x"b6",
          2687 => x"05",
          2688 => x"72",
          2689 => x"38",
          2690 => x"b6",
          2691 => x"05",
          2692 => x"39",
          2693 => x"08",
          2694 => x"70",
          2695 => x"08",
          2696 => x"29",
          2697 => x"08",
          2698 => x"70",
          2699 => x"a4",
          2700 => x"0c",
          2701 => x"08",
          2702 => x"70",
          2703 => x"71",
          2704 => x"51",
          2705 => x"53",
          2706 => x"b6",
          2707 => x"05",
          2708 => x"39",
          2709 => x"08",
          2710 => x"53",
          2711 => x"90",
          2712 => x"a4",
          2713 => x"08",
          2714 => x"a4",
          2715 => x"0c",
          2716 => x"08",
          2717 => x"82",
          2718 => x"fc",
          2719 => x"0c",
          2720 => x"82",
          2721 => x"ec",
          2722 => x"b6",
          2723 => x"05",
          2724 => x"98",
          2725 => x"0d",
          2726 => x"0c",
          2727 => x"0d",
          2728 => x"70",
          2729 => x"74",
          2730 => x"e3",
          2731 => x"75",
          2732 => x"d1",
          2733 => x"98",
          2734 => x"0c",
          2735 => x"54",
          2736 => x"74",
          2737 => x"a0",
          2738 => x"06",
          2739 => x"15",
          2740 => x"80",
          2741 => x"29",
          2742 => x"05",
          2743 => x"56",
          2744 => x"82",
          2745 => x"53",
          2746 => x"08",
          2747 => x"3f",
          2748 => x"08",
          2749 => x"16",
          2750 => x"81",
          2751 => x"38",
          2752 => x"81",
          2753 => x"54",
          2754 => x"c9",
          2755 => x"73",
          2756 => x"0c",
          2757 => x"04",
          2758 => x"73",
          2759 => x"26",
          2760 => x"71",
          2761 => x"95",
          2762 => x"71",
          2763 => x"9b",
          2764 => x"80",
          2765 => x"a4",
          2766 => x"39",
          2767 => x"51",
          2768 => x"82",
          2769 => x"80",
          2770 => x"9b",
          2771 => x"e4",
          2772 => x"e4",
          2773 => x"39",
          2774 => x"51",
          2775 => x"82",
          2776 => x"80",
          2777 => x"9c",
          2778 => x"c8",
          2779 => x"b8",
          2780 => x"39",
          2781 => x"51",
          2782 => x"9c",
          2783 => x"39",
          2784 => x"51",
          2785 => x"9d",
          2786 => x"39",
          2787 => x"51",
          2788 => x"9d",
          2789 => x"39",
          2790 => x"51",
          2791 => x"9e",
          2792 => x"39",
          2793 => x"51",
          2794 => x"9e",
          2795 => x"39",
          2796 => x"51",
          2797 => x"83",
          2798 => x"fb",
          2799 => x"79",
          2800 => x"87",
          2801 => x"38",
          2802 => x"87",
          2803 => x"90",
          2804 => x"52",
          2805 => x"ab",
          2806 => x"98",
          2807 => x"51",
          2808 => x"82",
          2809 => x"54",
          2810 => x"52",
          2811 => x"51",
          2812 => x"3f",
          2813 => x"04",
          2814 => x"66",
          2815 => x"80",
          2816 => x"5b",
          2817 => x"78",
          2818 => x"07",
          2819 => x"57",
          2820 => x"56",
          2821 => x"26",
          2822 => x"56",
          2823 => x"70",
          2824 => x"51",
          2825 => x"74",
          2826 => x"81",
          2827 => x"8c",
          2828 => x"56",
          2829 => x"3f",
          2830 => x"08",
          2831 => x"98",
          2832 => x"82",
          2833 => x"87",
          2834 => x"0c",
          2835 => x"08",
          2836 => x"d4",
          2837 => x"80",
          2838 => x"75",
          2839 => x"a3",
          2840 => x"98",
          2841 => x"b6",
          2842 => x"38",
          2843 => x"80",
          2844 => x"74",
          2845 => x"59",
          2846 => x"96",
          2847 => x"51",
          2848 => x"3f",
          2849 => x"78",
          2850 => x"7b",
          2851 => x"2a",
          2852 => x"57",
          2853 => x"80",
          2854 => x"82",
          2855 => x"87",
          2856 => x"08",
          2857 => x"fe",
          2858 => x"56",
          2859 => x"98",
          2860 => x"0d",
          2861 => x"0d",
          2862 => x"05",
          2863 => x"59",
          2864 => x"80",
          2865 => x"7b",
          2866 => x"3f",
          2867 => x"08",
          2868 => x"77",
          2869 => x"38",
          2870 => x"bf",
          2871 => x"82",
          2872 => x"82",
          2873 => x"82",
          2874 => x"82",
          2875 => x"54",
          2876 => x"08",
          2877 => x"e8",
          2878 => x"9e",
          2879 => x"b9",
          2880 => x"cd",
          2881 => x"55",
          2882 => x"b6",
          2883 => x"52",
          2884 => x"2d",
          2885 => x"08",
          2886 => x"79",
          2887 => x"b6",
          2888 => x"3d",
          2889 => x"3d",
          2890 => x"63",
          2891 => x"80",
          2892 => x"73",
          2893 => x"41",
          2894 => x"5e",
          2895 => x"52",
          2896 => x"51",
          2897 => x"3f",
          2898 => x"51",
          2899 => x"3f",
          2900 => x"79",
          2901 => x"38",
          2902 => x"89",
          2903 => x"2e",
          2904 => x"c6",
          2905 => x"53",
          2906 => x"8e",
          2907 => x"52",
          2908 => x"51",
          2909 => x"3f",
          2910 => x"9f",
          2911 => x"b8",
          2912 => x"15",
          2913 => x"39",
          2914 => x"72",
          2915 => x"38",
          2916 => x"82",
          2917 => x"ff",
          2918 => x"89",
          2919 => x"c0",
          2920 => x"b4",
          2921 => x"55",
          2922 => x"18",
          2923 => x"27",
          2924 => x"33",
          2925 => x"cc",
          2926 => x"9c",
          2927 => x"82",
          2928 => x"ff",
          2929 => x"81",
          2930 => x"cd",
          2931 => x"a0",
          2932 => x"3f",
          2933 => x"82",
          2934 => x"ff",
          2935 => x"80",
          2936 => x"27",
          2937 => x"74",
          2938 => x"55",
          2939 => x"72",
          2940 => x"38",
          2941 => x"53",
          2942 => x"83",
          2943 => x"75",
          2944 => x"81",
          2945 => x"53",
          2946 => x"90",
          2947 => x"fe",
          2948 => x"82",
          2949 => x"52",
          2950 => x"39",
          2951 => x"08",
          2952 => x"d7",
          2953 => x"15",
          2954 => x"39",
          2955 => x"51",
          2956 => x"78",
          2957 => x"5c",
          2958 => x"3f",
          2959 => x"08",
          2960 => x"98",
          2961 => x"76",
          2962 => x"81",
          2963 => x"9c",
          2964 => x"b6",
          2965 => x"2b",
          2966 => x"70",
          2967 => x"30",
          2968 => x"70",
          2969 => x"07",
          2970 => x"06",
          2971 => x"59",
          2972 => x"80",
          2973 => x"38",
          2974 => x"09",
          2975 => x"38",
          2976 => x"39",
          2977 => x"72",
          2978 => x"b2",
          2979 => x"72",
          2980 => x"0c",
          2981 => x"04",
          2982 => x"02",
          2983 => x"82",
          2984 => x"82",
          2985 => x"55",
          2986 => x"3f",
          2987 => x"22",
          2988 => x"3f",
          2989 => x"54",
          2990 => x"53",
          2991 => x"33",
          2992 => x"84",
          2993 => x"90",
          2994 => x"2e",
          2995 => x"d8",
          2996 => x"0d",
          2997 => x"0d",
          2998 => x"80",
          2999 => x"c0",
          3000 => x"98",
          3001 => x"a0",
          3002 => x"a3",
          3003 => x"98",
          3004 => x"81",
          3005 => x"06",
          3006 => x"80",
          3007 => x"81",
          3008 => x"3f",
          3009 => x"51",
          3010 => x"80",
          3011 => x"3f",
          3012 => x"70",
          3013 => x"52",
          3014 => x"92",
          3015 => x"97",
          3016 => x"a0",
          3017 => x"e7",
          3018 => x"97",
          3019 => x"83",
          3020 => x"06",
          3021 => x"80",
          3022 => x"81",
          3023 => x"3f",
          3024 => x"51",
          3025 => x"80",
          3026 => x"3f",
          3027 => x"70",
          3028 => x"52",
          3029 => x"92",
          3030 => x"97",
          3031 => x"a0",
          3032 => x"ab",
          3033 => x"97",
          3034 => x"85",
          3035 => x"06",
          3036 => x"80",
          3037 => x"81",
          3038 => x"3f",
          3039 => x"51",
          3040 => x"80",
          3041 => x"3f",
          3042 => x"70",
          3043 => x"52",
          3044 => x"92",
          3045 => x"96",
          3046 => x"a1",
          3047 => x"ef",
          3048 => x"96",
          3049 => x"87",
          3050 => x"06",
          3051 => x"80",
          3052 => x"81",
          3053 => x"3f",
          3054 => x"51",
          3055 => x"80",
          3056 => x"3f",
          3057 => x"70",
          3058 => x"52",
          3059 => x"92",
          3060 => x"96",
          3061 => x"a1",
          3062 => x"b3",
          3063 => x"96",
          3064 => x"c4",
          3065 => x"0d",
          3066 => x"0d",
          3067 => x"05",
          3068 => x"70",
          3069 => x"80",
          3070 => x"e2",
          3071 => x"0b",
          3072 => x"33",
          3073 => x"38",
          3074 => x"a1",
          3075 => x"cd",
          3076 => x"f8",
          3077 => x"b6",
          3078 => x"70",
          3079 => x"08",
          3080 => x"82",
          3081 => x"51",
          3082 => x"0b",
          3083 => x"34",
          3084 => x"b1",
          3085 => x"73",
          3086 => x"81",
          3087 => x"82",
          3088 => x"74",
          3089 => x"81",
          3090 => x"82",
          3091 => x"80",
          3092 => x"82",
          3093 => x"51",
          3094 => x"91",
          3095 => x"98",
          3096 => x"ab",
          3097 => x"0b",
          3098 => x"94",
          3099 => x"82",
          3100 => x"54",
          3101 => x"09",
          3102 => x"38",
          3103 => x"53",
          3104 => x"51",
          3105 => x"80",
          3106 => x"98",
          3107 => x"0d",
          3108 => x"0d",
          3109 => x"82",
          3110 => x"5f",
          3111 => x"7c",
          3112 => x"d5",
          3113 => x"98",
          3114 => x"06",
          3115 => x"2e",
          3116 => x"a3",
          3117 => x"59",
          3118 => x"a2",
          3119 => x"51",
          3120 => x"7c",
          3121 => x"82",
          3122 => x"80",
          3123 => x"82",
          3124 => x"7d",
          3125 => x"82",
          3126 => x"8d",
          3127 => x"70",
          3128 => x"a2",
          3129 => x"b1",
          3130 => x"3d",
          3131 => x"80",
          3132 => x"51",
          3133 => x"b4",
          3134 => x"05",
          3135 => x"3f",
          3136 => x"08",
          3137 => x"90",
          3138 => x"78",
          3139 => x"87",
          3140 => x"80",
          3141 => x"38",
          3142 => x"81",
          3143 => x"bd",
          3144 => x"78",
          3145 => x"ba",
          3146 => x"2e",
          3147 => x"8a",
          3148 => x"80",
          3149 => x"99",
          3150 => x"c0",
          3151 => x"38",
          3152 => x"82",
          3153 => x"bd",
          3154 => x"f9",
          3155 => x"38",
          3156 => x"24",
          3157 => x"80",
          3158 => x"88",
          3159 => x"f8",
          3160 => x"38",
          3161 => x"78",
          3162 => x"8a",
          3163 => x"81",
          3164 => x"38",
          3165 => x"2e",
          3166 => x"8a",
          3167 => x"81",
          3168 => x"fb",
          3169 => x"39",
          3170 => x"80",
          3171 => x"84",
          3172 => x"b8",
          3173 => x"98",
          3174 => x"fe",
          3175 => x"3d",
          3176 => x"53",
          3177 => x"51",
          3178 => x"82",
          3179 => x"80",
          3180 => x"38",
          3181 => x"f8",
          3182 => x"84",
          3183 => x"8c",
          3184 => x"98",
          3185 => x"82",
          3186 => x"42",
          3187 => x"51",
          3188 => x"3f",
          3189 => x"5a",
          3190 => x"81",
          3191 => x"59",
          3192 => x"84",
          3193 => x"7a",
          3194 => x"38",
          3195 => x"b4",
          3196 => x"11",
          3197 => x"05",
          3198 => x"3f",
          3199 => x"08",
          3200 => x"de",
          3201 => x"fe",
          3202 => x"ff",
          3203 => x"eb",
          3204 => x"b6",
          3205 => x"2e",
          3206 => x"b4",
          3207 => x"11",
          3208 => x"05",
          3209 => x"3f",
          3210 => x"08",
          3211 => x"b2",
          3212 => x"e0",
          3213 => x"a0",
          3214 => x"79",
          3215 => x"89",
          3216 => x"79",
          3217 => x"5b",
          3218 => x"61",
          3219 => x"eb",
          3220 => x"ff",
          3221 => x"ff",
          3222 => x"ea",
          3223 => x"b6",
          3224 => x"2e",
          3225 => x"b4",
          3226 => x"11",
          3227 => x"05",
          3228 => x"3f",
          3229 => x"08",
          3230 => x"e6",
          3231 => x"fe",
          3232 => x"ff",
          3233 => x"ea",
          3234 => x"b6",
          3235 => x"2e",
          3236 => x"82",
          3237 => x"ff",
          3238 => x"63",
          3239 => x"27",
          3240 => x"70",
          3241 => x"5e",
          3242 => x"7c",
          3243 => x"78",
          3244 => x"79",
          3245 => x"52",
          3246 => x"51",
          3247 => x"3f",
          3248 => x"81",
          3249 => x"d5",
          3250 => x"cd",
          3251 => x"92",
          3252 => x"ff",
          3253 => x"ff",
          3254 => x"e9",
          3255 => x"b6",
          3256 => x"df",
          3257 => x"84",
          3258 => x"80",
          3259 => x"82",
          3260 => x"44",
          3261 => x"82",
          3262 => x"59",
          3263 => x"88",
          3264 => x"c4",
          3265 => x"39",
          3266 => x"33",
          3267 => x"2e",
          3268 => x"b4",
          3269 => x"ab",
          3270 => x"87",
          3271 => x"80",
          3272 => x"82",
          3273 => x"44",
          3274 => x"b5",
          3275 => x"78",
          3276 => x"38",
          3277 => x"08",
          3278 => x"82",
          3279 => x"fc",
          3280 => x"b4",
          3281 => x"11",
          3282 => x"05",
          3283 => x"3f",
          3284 => x"08",
          3285 => x"82",
          3286 => x"59",
          3287 => x"89",
          3288 => x"c0",
          3289 => x"cc",
          3290 => x"85",
          3291 => x"80",
          3292 => x"82",
          3293 => x"43",
          3294 => x"b5",
          3295 => x"78",
          3296 => x"38",
          3297 => x"08",
          3298 => x"82",
          3299 => x"59",
          3300 => x"88",
          3301 => x"d8",
          3302 => x"39",
          3303 => x"33",
          3304 => x"2e",
          3305 => x"b4",
          3306 => x"88",
          3307 => x"ec",
          3308 => x"43",
          3309 => x"f8",
          3310 => x"84",
          3311 => x"8c",
          3312 => x"98",
          3313 => x"a7",
          3314 => x"5c",
          3315 => x"2e",
          3316 => x"5c",
          3317 => x"70",
          3318 => x"07",
          3319 => x"7f",
          3320 => x"5a",
          3321 => x"2e",
          3322 => x"a0",
          3323 => x"88",
          3324 => x"98",
          3325 => x"3f",
          3326 => x"54",
          3327 => x"52",
          3328 => x"a2",
          3329 => x"a4",
          3330 => x"39",
          3331 => x"80",
          3332 => x"84",
          3333 => x"b4",
          3334 => x"98",
          3335 => x"f9",
          3336 => x"3d",
          3337 => x"53",
          3338 => x"51",
          3339 => x"82",
          3340 => x"80",
          3341 => x"63",
          3342 => x"cb",
          3343 => x"34",
          3344 => x"44",
          3345 => x"fc",
          3346 => x"84",
          3347 => x"fc",
          3348 => x"98",
          3349 => x"f9",
          3350 => x"70",
          3351 => x"82",
          3352 => x"ff",
          3353 => x"82",
          3354 => x"53",
          3355 => x"79",
          3356 => x"b9",
          3357 => x"79",
          3358 => x"ae",
          3359 => x"38",
          3360 => x"9f",
          3361 => x"fe",
          3362 => x"ff",
          3363 => x"e6",
          3364 => x"b6",
          3365 => x"2e",
          3366 => x"59",
          3367 => x"05",
          3368 => x"63",
          3369 => x"ff",
          3370 => x"a3",
          3371 => x"b3",
          3372 => x"39",
          3373 => x"f4",
          3374 => x"84",
          3375 => x"bb",
          3376 => x"98",
          3377 => x"f8",
          3378 => x"3d",
          3379 => x"53",
          3380 => x"51",
          3381 => x"82",
          3382 => x"80",
          3383 => x"60",
          3384 => x"05",
          3385 => x"82",
          3386 => x"78",
          3387 => x"fe",
          3388 => x"ff",
          3389 => x"e0",
          3390 => x"b6",
          3391 => x"38",
          3392 => x"60",
          3393 => x"52",
          3394 => x"51",
          3395 => x"3f",
          3396 => x"08",
          3397 => x"52",
          3398 => x"aa",
          3399 => x"45",
          3400 => x"78",
          3401 => x"ba",
          3402 => x"26",
          3403 => x"82",
          3404 => x"39",
          3405 => x"f0",
          3406 => x"84",
          3407 => x"bb",
          3408 => x"98",
          3409 => x"92",
          3410 => x"02",
          3411 => x"79",
          3412 => x"5b",
          3413 => x"ff",
          3414 => x"a3",
          3415 => x"83",
          3416 => x"39",
          3417 => x"f4",
          3418 => x"84",
          3419 => x"8b",
          3420 => x"98",
          3421 => x"f6",
          3422 => x"3d",
          3423 => x"53",
          3424 => x"51",
          3425 => x"82",
          3426 => x"80",
          3427 => x"60",
          3428 => x"59",
          3429 => x"41",
          3430 => x"f0",
          3431 => x"84",
          3432 => x"d7",
          3433 => x"98",
          3434 => x"f6",
          3435 => x"70",
          3436 => x"82",
          3437 => x"ff",
          3438 => x"82",
          3439 => x"53",
          3440 => x"79",
          3441 => x"e5",
          3442 => x"79",
          3443 => x"ae",
          3444 => x"38",
          3445 => x"9b",
          3446 => x"fe",
          3447 => x"ff",
          3448 => x"de",
          3449 => x"b6",
          3450 => x"2e",
          3451 => x"60",
          3452 => x"60",
          3453 => x"ff",
          3454 => x"a3",
          3455 => x"e3",
          3456 => x"39",
          3457 => x"80",
          3458 => x"84",
          3459 => x"bc",
          3460 => x"98",
          3461 => x"f5",
          3462 => x"52",
          3463 => x"51",
          3464 => x"3f",
          3465 => x"04",
          3466 => x"80",
          3467 => x"84",
          3468 => x"98",
          3469 => x"98",
          3470 => x"f5",
          3471 => x"52",
          3472 => x"51",
          3473 => x"3f",
          3474 => x"2d",
          3475 => x"08",
          3476 => x"8e",
          3477 => x"98",
          3478 => x"a4",
          3479 => x"a6",
          3480 => x"fe",
          3481 => x"b0",
          3482 => x"3f",
          3483 => x"3f",
          3484 => x"82",
          3485 => x"c2",
          3486 => x"59",
          3487 => x"91",
          3488 => x"de",
          3489 => x"79",
          3490 => x"80",
          3491 => x"38",
          3492 => x"59",
          3493 => x"81",
          3494 => x"3d",
          3495 => x"51",
          3496 => x"82",
          3497 => x"5c",
          3498 => x"82",
          3499 => x"7a",
          3500 => x"38",
          3501 => x"8c",
          3502 => x"39",
          3503 => x"ad",
          3504 => x"39",
          3505 => x"56",
          3506 => x"a4",
          3507 => x"53",
          3508 => x"52",
          3509 => x"b0",
          3510 => x"a8",
          3511 => x"39",
          3512 => x"3d",
          3513 => x"51",
          3514 => x"ab",
          3515 => x"82",
          3516 => x"80",
          3517 => x"f8",
          3518 => x"ff",
          3519 => x"ff",
          3520 => x"93",
          3521 => x"80",
          3522 => x"84",
          3523 => x"ff",
          3524 => x"ff",
          3525 => x"82",
          3526 => x"82",
          3527 => x"80",
          3528 => x"80",
          3529 => x"80",
          3530 => x"80",
          3531 => x"ff",
          3532 => x"eb",
          3533 => x"b6",
          3534 => x"b6",
          3535 => x"70",
          3536 => x"07",
          3537 => x"5b",
          3538 => x"5a",
          3539 => x"83",
          3540 => x"78",
          3541 => x"78",
          3542 => x"38",
          3543 => x"81",
          3544 => x"59",
          3545 => x"38",
          3546 => x"7d",
          3547 => x"59",
          3548 => x"7e",
          3549 => x"81",
          3550 => x"38",
          3551 => x"51",
          3552 => x"f2",
          3553 => x"3d",
          3554 => x"82",
          3555 => x"87",
          3556 => x"70",
          3557 => x"87",
          3558 => x"72",
          3559 => x"3f",
          3560 => x"08",
          3561 => x"08",
          3562 => x"84",
          3563 => x"51",
          3564 => x"72",
          3565 => x"08",
          3566 => x"87",
          3567 => x"70",
          3568 => x"87",
          3569 => x"72",
          3570 => x"3f",
          3571 => x"08",
          3572 => x"08",
          3573 => x"84",
          3574 => x"51",
          3575 => x"72",
          3576 => x"08",
          3577 => x"8c",
          3578 => x"87",
          3579 => x"0c",
          3580 => x"0b",
          3581 => x"94",
          3582 => x"8b",
          3583 => x"f7",
          3584 => x"84",
          3585 => x"34",
          3586 => x"cd",
          3587 => x"3d",
          3588 => x"0c",
          3589 => x"82",
          3590 => x"54",
          3591 => x"92",
          3592 => x"a5",
          3593 => x"bf",
          3594 => x"a5",
          3595 => x"bf",
          3596 => x"dd",
          3597 => x"e3",
          3598 => x"ec",
          3599 => x"d1",
          3600 => x"fe",
          3601 => x"52",
          3602 => x"88",
          3603 => x"d8",
          3604 => x"98",
          3605 => x"06",
          3606 => x"14",
          3607 => x"80",
          3608 => x"71",
          3609 => x"0c",
          3610 => x"04",
          3611 => x"76",
          3612 => x"55",
          3613 => x"54",
          3614 => x"81",
          3615 => x"33",
          3616 => x"2e",
          3617 => x"86",
          3618 => x"53",
          3619 => x"33",
          3620 => x"2e",
          3621 => x"86",
          3622 => x"53",
          3623 => x"52",
          3624 => x"09",
          3625 => x"38",
          3626 => x"12",
          3627 => x"33",
          3628 => x"a2",
          3629 => x"81",
          3630 => x"2e",
          3631 => x"ea",
          3632 => x"81",
          3633 => x"72",
          3634 => x"70",
          3635 => x"38",
          3636 => x"80",
          3637 => x"73",
          3638 => x"72",
          3639 => x"70",
          3640 => x"81",
          3641 => x"81",
          3642 => x"32",
          3643 => x"80",
          3644 => x"51",
          3645 => x"80",
          3646 => x"80",
          3647 => x"05",
          3648 => x"75",
          3649 => x"70",
          3650 => x"0c",
          3651 => x"04",
          3652 => x"76",
          3653 => x"80",
          3654 => x"86",
          3655 => x"52",
          3656 => x"d7",
          3657 => x"98",
          3658 => x"80",
          3659 => x"74",
          3660 => x"b6",
          3661 => x"3d",
          3662 => x"3d",
          3663 => x"11",
          3664 => x"52",
          3665 => x"70",
          3666 => x"98",
          3667 => x"33",
          3668 => x"82",
          3669 => x"26",
          3670 => x"84",
          3671 => x"83",
          3672 => x"26",
          3673 => x"85",
          3674 => x"84",
          3675 => x"26",
          3676 => x"86",
          3677 => x"85",
          3678 => x"26",
          3679 => x"88",
          3680 => x"86",
          3681 => x"e7",
          3682 => x"38",
          3683 => x"54",
          3684 => x"87",
          3685 => x"cc",
          3686 => x"87",
          3687 => x"0c",
          3688 => x"c0",
          3689 => x"82",
          3690 => x"c0",
          3691 => x"83",
          3692 => x"c0",
          3693 => x"84",
          3694 => x"c0",
          3695 => x"85",
          3696 => x"c0",
          3697 => x"86",
          3698 => x"c0",
          3699 => x"74",
          3700 => x"a4",
          3701 => x"c0",
          3702 => x"80",
          3703 => x"98",
          3704 => x"52",
          3705 => x"98",
          3706 => x"0d",
          3707 => x"0d",
          3708 => x"c0",
          3709 => x"81",
          3710 => x"c0",
          3711 => x"5e",
          3712 => x"87",
          3713 => x"08",
          3714 => x"1c",
          3715 => x"98",
          3716 => x"79",
          3717 => x"87",
          3718 => x"08",
          3719 => x"1c",
          3720 => x"98",
          3721 => x"79",
          3722 => x"87",
          3723 => x"08",
          3724 => x"1c",
          3725 => x"98",
          3726 => x"7b",
          3727 => x"87",
          3728 => x"08",
          3729 => x"1c",
          3730 => x"0c",
          3731 => x"ff",
          3732 => x"83",
          3733 => x"58",
          3734 => x"57",
          3735 => x"56",
          3736 => x"55",
          3737 => x"54",
          3738 => x"53",
          3739 => x"ff",
          3740 => x"a5",
          3741 => x"9e",
          3742 => x"3d",
          3743 => x"3d",
          3744 => x"05",
          3745 => x"b8",
          3746 => x"ff",
          3747 => x"55",
          3748 => x"84",
          3749 => x"2e",
          3750 => x"c0",
          3751 => x"70",
          3752 => x"2a",
          3753 => x"53",
          3754 => x"80",
          3755 => x"71",
          3756 => x"81",
          3757 => x"70",
          3758 => x"81",
          3759 => x"06",
          3760 => x"80",
          3761 => x"71",
          3762 => x"81",
          3763 => x"70",
          3764 => x"73",
          3765 => x"51",
          3766 => x"80",
          3767 => x"2e",
          3768 => x"c0",
          3769 => x"74",
          3770 => x"82",
          3771 => x"87",
          3772 => x"ff",
          3773 => x"8f",
          3774 => x"30",
          3775 => x"51",
          3776 => x"82",
          3777 => x"83",
          3778 => x"f9",
          3779 => x"a7",
          3780 => x"77",
          3781 => x"81",
          3782 => x"7a",
          3783 => x"eb",
          3784 => x"b8",
          3785 => x"ff",
          3786 => x"87",
          3787 => x"53",
          3788 => x"86",
          3789 => x"94",
          3790 => x"08",
          3791 => x"70",
          3792 => x"56",
          3793 => x"2e",
          3794 => x"91",
          3795 => x"06",
          3796 => x"d7",
          3797 => x"32",
          3798 => x"51",
          3799 => x"2e",
          3800 => x"93",
          3801 => x"06",
          3802 => x"ff",
          3803 => x"81",
          3804 => x"87",
          3805 => x"54",
          3806 => x"86",
          3807 => x"94",
          3808 => x"74",
          3809 => x"82",
          3810 => x"89",
          3811 => x"f9",
          3812 => x"54",
          3813 => x"70",
          3814 => x"53",
          3815 => x"77",
          3816 => x"38",
          3817 => x"06",
          3818 => x"b4",
          3819 => x"81",
          3820 => x"57",
          3821 => x"c0",
          3822 => x"75",
          3823 => x"38",
          3824 => x"94",
          3825 => x"70",
          3826 => x"81",
          3827 => x"52",
          3828 => x"8c",
          3829 => x"2a",
          3830 => x"51",
          3831 => x"38",
          3832 => x"70",
          3833 => x"51",
          3834 => x"8d",
          3835 => x"2a",
          3836 => x"51",
          3837 => x"be",
          3838 => x"ff",
          3839 => x"c0",
          3840 => x"70",
          3841 => x"38",
          3842 => x"90",
          3843 => x"0c",
          3844 => x"33",
          3845 => x"06",
          3846 => x"70",
          3847 => x"76",
          3848 => x"0c",
          3849 => x"04",
          3850 => x"82",
          3851 => x"70",
          3852 => x"54",
          3853 => x"94",
          3854 => x"80",
          3855 => x"87",
          3856 => x"51",
          3857 => x"82",
          3858 => x"06",
          3859 => x"70",
          3860 => x"38",
          3861 => x"06",
          3862 => x"94",
          3863 => x"80",
          3864 => x"87",
          3865 => x"52",
          3866 => x"81",
          3867 => x"b6",
          3868 => x"84",
          3869 => x"ff",
          3870 => x"b6",
          3871 => x"ff",
          3872 => x"98",
          3873 => x"3d",
          3874 => x"b8",
          3875 => x"ff",
          3876 => x"87",
          3877 => x"52",
          3878 => x"86",
          3879 => x"94",
          3880 => x"08",
          3881 => x"70",
          3882 => x"51",
          3883 => x"70",
          3884 => x"38",
          3885 => x"06",
          3886 => x"94",
          3887 => x"80",
          3888 => x"87",
          3889 => x"52",
          3890 => x"98",
          3891 => x"2c",
          3892 => x"71",
          3893 => x"0c",
          3894 => x"04",
          3895 => x"87",
          3896 => x"08",
          3897 => x"8a",
          3898 => x"70",
          3899 => x"b4",
          3900 => x"9e",
          3901 => x"b4",
          3902 => x"c0",
          3903 => x"82",
          3904 => x"87",
          3905 => x"08",
          3906 => x"0c",
          3907 => x"98",
          3908 => x"c8",
          3909 => x"9e",
          3910 => x"b4",
          3911 => x"c0",
          3912 => x"82",
          3913 => x"87",
          3914 => x"08",
          3915 => x"0c",
          3916 => x"b0",
          3917 => x"d8",
          3918 => x"9e",
          3919 => x"b4",
          3920 => x"c0",
          3921 => x"82",
          3922 => x"87",
          3923 => x"08",
          3924 => x"0c",
          3925 => x"c0",
          3926 => x"e8",
          3927 => x"9e",
          3928 => x"b4",
          3929 => x"c0",
          3930 => x"51",
          3931 => x"f0",
          3932 => x"9e",
          3933 => x"b4",
          3934 => x"c0",
          3935 => x"82",
          3936 => x"87",
          3937 => x"08",
          3938 => x"0c",
          3939 => x"b5",
          3940 => x"0b",
          3941 => x"90",
          3942 => x"80",
          3943 => x"52",
          3944 => x"2e",
          3945 => x"52",
          3946 => x"81",
          3947 => x"87",
          3948 => x"08",
          3949 => x"0a",
          3950 => x"52",
          3951 => x"83",
          3952 => x"71",
          3953 => x"34",
          3954 => x"c0",
          3955 => x"70",
          3956 => x"06",
          3957 => x"70",
          3958 => x"38",
          3959 => x"82",
          3960 => x"80",
          3961 => x"9e",
          3962 => x"88",
          3963 => x"51",
          3964 => x"80",
          3965 => x"81",
          3966 => x"b5",
          3967 => x"0b",
          3968 => x"90",
          3969 => x"80",
          3970 => x"52",
          3971 => x"2e",
          3972 => x"52",
          3973 => x"85",
          3974 => x"87",
          3975 => x"08",
          3976 => x"80",
          3977 => x"52",
          3978 => x"83",
          3979 => x"71",
          3980 => x"34",
          3981 => x"c0",
          3982 => x"70",
          3983 => x"06",
          3984 => x"70",
          3985 => x"38",
          3986 => x"82",
          3987 => x"80",
          3988 => x"9e",
          3989 => x"82",
          3990 => x"51",
          3991 => x"80",
          3992 => x"81",
          3993 => x"b5",
          3994 => x"0b",
          3995 => x"90",
          3996 => x"80",
          3997 => x"52",
          3998 => x"2e",
          3999 => x"52",
          4000 => x"89",
          4001 => x"87",
          4002 => x"08",
          4003 => x"80",
          4004 => x"52",
          4005 => x"83",
          4006 => x"71",
          4007 => x"34",
          4008 => x"c0",
          4009 => x"70",
          4010 => x"51",
          4011 => x"80",
          4012 => x"81",
          4013 => x"b5",
          4014 => x"c0",
          4015 => x"70",
          4016 => x"70",
          4017 => x"51",
          4018 => x"b5",
          4019 => x"0b",
          4020 => x"90",
          4021 => x"80",
          4022 => x"52",
          4023 => x"83",
          4024 => x"71",
          4025 => x"34",
          4026 => x"90",
          4027 => x"f0",
          4028 => x"2a",
          4029 => x"70",
          4030 => x"34",
          4031 => x"c0",
          4032 => x"70",
          4033 => x"52",
          4034 => x"2e",
          4035 => x"52",
          4036 => x"8f",
          4037 => x"9e",
          4038 => x"87",
          4039 => x"70",
          4040 => x"34",
          4041 => x"04",
          4042 => x"82",
          4043 => x"ff",
          4044 => x"82",
          4045 => x"54",
          4046 => x"89",
          4047 => x"ec",
          4048 => x"94",
          4049 => x"80",
          4050 => x"97",
          4051 => x"82",
          4052 => x"80",
          4053 => x"82",
          4054 => x"82",
          4055 => x"11",
          4056 => x"a6",
          4057 => x"94",
          4058 => x"b5",
          4059 => x"73",
          4060 => x"38",
          4061 => x"08",
          4062 => x"08",
          4063 => x"82",
          4064 => x"ff",
          4065 => x"82",
          4066 => x"54",
          4067 => x"94",
          4068 => x"bc",
          4069 => x"c0",
          4070 => x"52",
          4071 => x"51",
          4072 => x"3f",
          4073 => x"33",
          4074 => x"2e",
          4075 => x"b4",
          4076 => x"b4",
          4077 => x"54",
          4078 => x"ec",
          4079 => x"98",
          4080 => x"86",
          4081 => x"80",
          4082 => x"82",
          4083 => x"82",
          4084 => x"11",
          4085 => x"a7",
          4086 => x"93",
          4087 => x"b5",
          4088 => x"73",
          4089 => x"38",
          4090 => x"33",
          4091 => x"a4",
          4092 => x"e4",
          4093 => x"8f",
          4094 => x"80",
          4095 => x"82",
          4096 => x"52",
          4097 => x"51",
          4098 => x"3f",
          4099 => x"33",
          4100 => x"2e",
          4101 => x"b5",
          4102 => x"82",
          4103 => x"ff",
          4104 => x"82",
          4105 => x"54",
          4106 => x"89",
          4107 => x"84",
          4108 => x"af",
          4109 => x"83",
          4110 => x"80",
          4111 => x"82",
          4112 => x"ff",
          4113 => x"82",
          4114 => x"54",
          4115 => x"89",
          4116 => x"a4",
          4117 => x"8b",
          4118 => x"89",
          4119 => x"80",
          4120 => x"82",
          4121 => x"ff",
          4122 => x"82",
          4123 => x"54",
          4124 => x"89",
          4125 => x"b8",
          4126 => x"e7",
          4127 => x"c0",
          4128 => x"df",
          4129 => x"e4",
          4130 => x"a8",
          4131 => x"92",
          4132 => x"b4",
          4133 => x"82",
          4134 => x"ff",
          4135 => x"82",
          4136 => x"52",
          4137 => x"51",
          4138 => x"3f",
          4139 => x"51",
          4140 => x"3f",
          4141 => x"22",
          4142 => x"cc",
          4143 => x"98",
          4144 => x"f4",
          4145 => x"84",
          4146 => x"51",
          4147 => x"82",
          4148 => x"bd",
          4149 => x"76",
          4150 => x"54",
          4151 => x"08",
          4152 => x"f4",
          4153 => x"f0",
          4154 => x"87",
          4155 => x"80",
          4156 => x"82",
          4157 => x"56",
          4158 => x"52",
          4159 => x"83",
          4160 => x"98",
          4161 => x"c0",
          4162 => x"31",
          4163 => x"b6",
          4164 => x"82",
          4165 => x"ff",
          4166 => x"82",
          4167 => x"54",
          4168 => x"a9",
          4169 => x"fc",
          4170 => x"84",
          4171 => x"51",
          4172 => x"82",
          4173 => x"bd",
          4174 => x"76",
          4175 => x"54",
          4176 => x"08",
          4177 => x"cc",
          4178 => x"8c",
          4179 => x"ff",
          4180 => x"87",
          4181 => x"fe",
          4182 => x"92",
          4183 => x"05",
          4184 => x"26",
          4185 => x"84",
          4186 => x"9c",
          4187 => x"08",
          4188 => x"f8",
          4189 => x"82",
          4190 => x"97",
          4191 => x"88",
          4192 => x"82",
          4193 => x"8b",
          4194 => x"94",
          4195 => x"82",
          4196 => x"ff",
          4197 => x"84",
          4198 => x"71",
          4199 => x"04",
          4200 => x"c0",
          4201 => x"04",
          4202 => x"08",
          4203 => x"84",
          4204 => x"3d",
          4205 => x"2b",
          4206 => x"79",
          4207 => x"98",
          4208 => x"13",
          4209 => x"51",
          4210 => x"51",
          4211 => x"82",
          4212 => x"33",
          4213 => x"74",
          4214 => x"82",
          4215 => x"08",
          4216 => x"05",
          4217 => x"71",
          4218 => x"52",
          4219 => x"09",
          4220 => x"38",
          4221 => x"82",
          4222 => x"85",
          4223 => x"fb",
          4224 => x"02",
          4225 => x"05",
          4226 => x"55",
          4227 => x"80",
          4228 => x"82",
          4229 => x"52",
          4230 => x"af",
          4231 => x"cd",
          4232 => x"a0",
          4233 => x"8a",
          4234 => x"ec",
          4235 => x"51",
          4236 => x"3f",
          4237 => x"05",
          4238 => x"34",
          4239 => x"06",
          4240 => x"77",
          4241 => x"90",
          4242 => x"34",
          4243 => x"04",
          4244 => x"7c",
          4245 => x"b7",
          4246 => x"88",
          4247 => x"33",
          4248 => x"33",
          4249 => x"82",
          4250 => x"70",
          4251 => x"59",
          4252 => x"74",
          4253 => x"38",
          4254 => x"fa",
          4255 => x"f0",
          4256 => x"29",
          4257 => x"05",
          4258 => x"54",
          4259 => x"9d",
          4260 => x"b6",
          4261 => x"0c",
          4262 => x"33",
          4263 => x"82",
          4264 => x"70",
          4265 => x"5a",
          4266 => x"a7",
          4267 => x"78",
          4268 => x"ff",
          4269 => x"82",
          4270 => x"81",
          4271 => x"82",
          4272 => x"74",
          4273 => x"55",
          4274 => x"87",
          4275 => x"82",
          4276 => x"77",
          4277 => x"38",
          4278 => x"08",
          4279 => x"2e",
          4280 => x"b5",
          4281 => x"74",
          4282 => x"3d",
          4283 => x"76",
          4284 => x"75",
          4285 => x"88",
          4286 => x"ec",
          4287 => x"51",
          4288 => x"3f",
          4289 => x"08",
          4290 => x"e5",
          4291 => x"0d",
          4292 => x"0d",
          4293 => x"53",
          4294 => x"08",
          4295 => x"2e",
          4296 => x"51",
          4297 => x"80",
          4298 => x"14",
          4299 => x"54",
          4300 => x"e6",
          4301 => x"82",
          4302 => x"82",
          4303 => x"52",
          4304 => x"95",
          4305 => x"80",
          4306 => x"82",
          4307 => x"51",
          4308 => x"80",
          4309 => x"ec",
          4310 => x"0d",
          4311 => x"0d",
          4312 => x"52",
          4313 => x"08",
          4314 => x"b2",
          4315 => x"98",
          4316 => x"38",
          4317 => x"08",
          4318 => x"52",
          4319 => x"52",
          4320 => x"80",
          4321 => x"98",
          4322 => x"ba",
          4323 => x"ff",
          4324 => x"82",
          4325 => x"55",
          4326 => x"b6",
          4327 => x"9d",
          4328 => x"98",
          4329 => x"70",
          4330 => x"80",
          4331 => x"53",
          4332 => x"17",
          4333 => x"52",
          4334 => x"9c",
          4335 => x"2e",
          4336 => x"ff",
          4337 => x"3d",
          4338 => x"3d",
          4339 => x"08",
          4340 => x"5a",
          4341 => x"58",
          4342 => x"82",
          4343 => x"51",
          4344 => x"3f",
          4345 => x"08",
          4346 => x"ff",
          4347 => x"ec",
          4348 => x"80",
          4349 => x"3d",
          4350 => x"81",
          4351 => x"82",
          4352 => x"80",
          4353 => x"75",
          4354 => x"f9",
          4355 => x"98",
          4356 => x"58",
          4357 => x"82",
          4358 => x"25",
          4359 => x"b6",
          4360 => x"05",
          4361 => x"55",
          4362 => x"74",
          4363 => x"70",
          4364 => x"2a",
          4365 => x"78",
          4366 => x"38",
          4367 => x"38",
          4368 => x"08",
          4369 => x"53",
          4370 => x"d2",
          4371 => x"98",
          4372 => x"89",
          4373 => x"a4",
          4374 => x"fc",
          4375 => x"2e",
          4376 => x"9b",
          4377 => x"79",
          4378 => x"87",
          4379 => x"ff",
          4380 => x"ab",
          4381 => x"82",
          4382 => x"74",
          4383 => x"77",
          4384 => x"0c",
          4385 => x"04",
          4386 => x"7c",
          4387 => x"71",
          4388 => x"59",
          4389 => x"a0",
          4390 => x"06",
          4391 => x"33",
          4392 => x"77",
          4393 => x"38",
          4394 => x"5b",
          4395 => x"56",
          4396 => x"a0",
          4397 => x"06",
          4398 => x"75",
          4399 => x"80",
          4400 => x"29",
          4401 => x"05",
          4402 => x"55",
          4403 => x"3f",
          4404 => x"08",
          4405 => x"74",
          4406 => x"b5",
          4407 => x"b6",
          4408 => x"c5",
          4409 => x"33",
          4410 => x"2e",
          4411 => x"82",
          4412 => x"b5",
          4413 => x"3f",
          4414 => x"1a",
          4415 => x"fc",
          4416 => x"05",
          4417 => x"3f",
          4418 => x"08",
          4419 => x"38",
          4420 => x"78",
          4421 => x"fd",
          4422 => x"b6",
          4423 => x"ff",
          4424 => x"85",
          4425 => x"91",
          4426 => x"70",
          4427 => x"51",
          4428 => x"27",
          4429 => x"80",
          4430 => x"b6",
          4431 => x"3d",
          4432 => x"3d",
          4433 => x"08",
          4434 => x"b4",
          4435 => x"5f",
          4436 => x"af",
          4437 => x"b5",
          4438 => x"b5",
          4439 => x"5b",
          4440 => x"38",
          4441 => x"e8",
          4442 => x"73",
          4443 => x"55",
          4444 => x"81",
          4445 => x"70",
          4446 => x"56",
          4447 => x"81",
          4448 => x"51",
          4449 => x"82",
          4450 => x"82",
          4451 => x"82",
          4452 => x"80",
          4453 => x"38",
          4454 => x"52",
          4455 => x"08",
          4456 => x"fa",
          4457 => x"98",
          4458 => x"8c",
          4459 => x"d0",
          4460 => x"af",
          4461 => x"39",
          4462 => x"08",
          4463 => x"ec",
          4464 => x"f8",
          4465 => x"70",
          4466 => x"87",
          4467 => x"b6",
          4468 => x"82",
          4469 => x"74",
          4470 => x"06",
          4471 => x"82",
          4472 => x"51",
          4473 => x"3f",
          4474 => x"08",
          4475 => x"82",
          4476 => x"25",
          4477 => x"b6",
          4478 => x"05",
          4479 => x"55",
          4480 => x"80",
          4481 => x"ff",
          4482 => x"51",
          4483 => x"81",
          4484 => x"ff",
          4485 => x"93",
          4486 => x"38",
          4487 => x"ff",
          4488 => x"06",
          4489 => x"86",
          4490 => x"b5",
          4491 => x"8c",
          4492 => x"ec",
          4493 => x"84",
          4494 => x"3f",
          4495 => x"ec",
          4496 => x"b6",
          4497 => x"2b",
          4498 => x"51",
          4499 => x"2e",
          4500 => x"81",
          4501 => x"cd",
          4502 => x"98",
          4503 => x"2c",
          4504 => x"33",
          4505 => x"70",
          4506 => x"98",
          4507 => x"84",
          4508 => x"a4",
          4509 => x"15",
          4510 => x"51",
          4511 => x"59",
          4512 => x"58",
          4513 => x"78",
          4514 => x"38",
          4515 => x"b4",
          4516 => x"80",
          4517 => x"ff",
          4518 => x"98",
          4519 => x"80",
          4520 => x"ce",
          4521 => x"74",
          4522 => x"f6",
          4523 => x"b6",
          4524 => x"ff",
          4525 => x"80",
          4526 => x"74",
          4527 => x"34",
          4528 => x"39",
          4529 => x"0a",
          4530 => x"0a",
          4531 => x"2c",
          4532 => x"06",
          4533 => x"73",
          4534 => x"38",
          4535 => x"52",
          4536 => x"ce",
          4537 => x"98",
          4538 => x"06",
          4539 => x"38",
          4540 => x"56",
          4541 => x"80",
          4542 => x"1c",
          4543 => x"cd",
          4544 => x"98",
          4545 => x"2c",
          4546 => x"33",
          4547 => x"70",
          4548 => x"10",
          4549 => x"2b",
          4550 => x"11",
          4551 => x"51",
          4552 => x"51",
          4553 => x"2e",
          4554 => x"fe",
          4555 => x"ab",
          4556 => x"7d",
          4557 => x"82",
          4558 => x"80",
          4559 => x"c0",
          4560 => x"75",
          4561 => x"34",
          4562 => x"c0",
          4563 => x"3d",
          4564 => x"0c",
          4565 => x"95",
          4566 => x"38",
          4567 => x"82",
          4568 => x"54",
          4569 => x"82",
          4570 => x"54",
          4571 => x"fd",
          4572 => x"cd",
          4573 => x"73",
          4574 => x"38",
          4575 => x"70",
          4576 => x"55",
          4577 => x"9e",
          4578 => x"54",
          4579 => x"15",
          4580 => x"80",
          4581 => x"ff",
          4582 => x"98",
          4583 => x"cc",
          4584 => x"55",
          4585 => x"cd",
          4586 => x"11",
          4587 => x"82",
          4588 => x"73",
          4589 => x"3d",
          4590 => x"82",
          4591 => x"54",
          4592 => x"89",
          4593 => x"54",
          4594 => x"c8",
          4595 => x"cc",
          4596 => x"80",
          4597 => x"ff",
          4598 => x"98",
          4599 => x"c8",
          4600 => x"56",
          4601 => x"25",
          4602 => x"cd",
          4603 => x"74",
          4604 => x"52",
          4605 => x"ba",
          4606 => x"80",
          4607 => x"80",
          4608 => x"98",
          4609 => x"c8",
          4610 => x"55",
          4611 => x"da",
          4612 => x"cc",
          4613 => x"2b",
          4614 => x"82",
          4615 => x"5a",
          4616 => x"74",
          4617 => x"94",
          4618 => x"ec",
          4619 => x"51",
          4620 => x"3f",
          4621 => x"0a",
          4622 => x"0a",
          4623 => x"2c",
          4624 => x"33",
          4625 => x"73",
          4626 => x"38",
          4627 => x"83",
          4628 => x"0b",
          4629 => x"82",
          4630 => x"80",
          4631 => x"ec",
          4632 => x"3f",
          4633 => x"82",
          4634 => x"70",
          4635 => x"55",
          4636 => x"2e",
          4637 => x"82",
          4638 => x"ff",
          4639 => x"82",
          4640 => x"ff",
          4641 => x"82",
          4642 => x"82",
          4643 => x"52",
          4644 => x"a2",
          4645 => x"cd",
          4646 => x"98",
          4647 => x"2c",
          4648 => x"33",
          4649 => x"57",
          4650 => x"ad",
          4651 => x"54",
          4652 => x"74",
          4653 => x"ec",
          4654 => x"33",
          4655 => x"f2",
          4656 => x"80",
          4657 => x"80",
          4658 => x"98",
          4659 => x"c8",
          4660 => x"55",
          4661 => x"d5",
          4662 => x"ec",
          4663 => x"51",
          4664 => x"3f",
          4665 => x"33",
          4666 => x"70",
          4667 => x"cd",
          4668 => x"51",
          4669 => x"74",
          4670 => x"38",
          4671 => x"08",
          4672 => x"ff",
          4673 => x"74",
          4674 => x"29",
          4675 => x"05",
          4676 => x"82",
          4677 => x"58",
          4678 => x"75",
          4679 => x"fa",
          4680 => x"cd",
          4681 => x"05",
          4682 => x"34",
          4683 => x"08",
          4684 => x"ff",
          4685 => x"82",
          4686 => x"79",
          4687 => x"3f",
          4688 => x"08",
          4689 => x"54",
          4690 => x"82",
          4691 => x"54",
          4692 => x"8f",
          4693 => x"73",
          4694 => x"f1",
          4695 => x"39",
          4696 => x"80",
          4697 => x"cc",
          4698 => x"82",
          4699 => x"79",
          4700 => x"0c",
          4701 => x"04",
          4702 => x"33",
          4703 => x"2e",
          4704 => x"82",
          4705 => x"52",
          4706 => x"a0",
          4707 => x"cd",
          4708 => x"05",
          4709 => x"cd",
          4710 => x"81",
          4711 => x"dd",
          4712 => x"cc",
          4713 => x"c8",
          4714 => x"73",
          4715 => x"8c",
          4716 => x"54",
          4717 => x"c8",
          4718 => x"2b",
          4719 => x"75",
          4720 => x"56",
          4721 => x"74",
          4722 => x"74",
          4723 => x"14",
          4724 => x"82",
          4725 => x"52",
          4726 => x"ff",
          4727 => x"74",
          4728 => x"29",
          4729 => x"05",
          4730 => x"82",
          4731 => x"58",
          4732 => x"75",
          4733 => x"82",
          4734 => x"52",
          4735 => x"9f",
          4736 => x"cd",
          4737 => x"98",
          4738 => x"2c",
          4739 => x"33",
          4740 => x"57",
          4741 => x"f8",
          4742 => x"cd",
          4743 => x"88",
          4744 => x"8e",
          4745 => x"80",
          4746 => x"80",
          4747 => x"98",
          4748 => x"c8",
          4749 => x"55",
          4750 => x"de",
          4751 => x"39",
          4752 => x"33",
          4753 => x"06",
          4754 => x"33",
          4755 => x"74",
          4756 => x"e8",
          4757 => x"ec",
          4758 => x"14",
          4759 => x"cd",
          4760 => x"1a",
          4761 => x"54",
          4762 => x"3f",
          4763 => x"33",
          4764 => x"06",
          4765 => x"33",
          4766 => x"75",
          4767 => x"38",
          4768 => x"82",
          4769 => x"80",
          4770 => x"ec",
          4771 => x"3f",
          4772 => x"cd",
          4773 => x"0b",
          4774 => x"34",
          4775 => x"7a",
          4776 => x"b5",
          4777 => x"74",
          4778 => x"38",
          4779 => x"a6",
          4780 => x"b6",
          4781 => x"cd",
          4782 => x"b6",
          4783 => x"ff",
          4784 => x"53",
          4785 => x"51",
          4786 => x"3f",
          4787 => x"c0",
          4788 => x"29",
          4789 => x"05",
          4790 => x"56",
          4791 => x"2e",
          4792 => x"51",
          4793 => x"3f",
          4794 => x"08",
          4795 => x"34",
          4796 => x"08",
          4797 => x"81",
          4798 => x"52",
          4799 => x"a7",
          4800 => x"1b",
          4801 => x"39",
          4802 => x"74",
          4803 => x"ac",
          4804 => x"ff",
          4805 => x"99",
          4806 => x"2e",
          4807 => x"ae",
          4808 => x"98",
          4809 => x"80",
          4810 => x"74",
          4811 => x"d5",
          4812 => x"98",
          4813 => x"c8",
          4814 => x"98",
          4815 => x"06",
          4816 => x"74",
          4817 => x"ff",
          4818 => x"80",
          4819 => x"84",
          4820 => x"9c",
          4821 => x"56",
          4822 => x"2e",
          4823 => x"51",
          4824 => x"3f",
          4825 => x"08",
          4826 => x"34",
          4827 => x"08",
          4828 => x"81",
          4829 => x"52",
          4830 => x"a6",
          4831 => x"1b",
          4832 => x"ff",
          4833 => x"39",
          4834 => x"c8",
          4835 => x"34",
          4836 => x"53",
          4837 => x"33",
          4838 => x"ec",
          4839 => x"9c",
          4840 => x"cc",
          4841 => x"ff",
          4842 => x"c8",
          4843 => x"54",
          4844 => x"f5",
          4845 => x"cd",
          4846 => x"81",
          4847 => x"82",
          4848 => x"74",
          4849 => x"52",
          4850 => x"e6",
          4851 => x"39",
          4852 => x"33",
          4853 => x"2e",
          4854 => x"82",
          4855 => x"52",
          4856 => x"9b",
          4857 => x"cd",
          4858 => x"05",
          4859 => x"cd",
          4860 => x"c8",
          4861 => x"0d",
          4862 => x"0b",
          4863 => x"0c",
          4864 => x"82",
          4865 => x"a0",
          4866 => x"52",
          4867 => x"51",
          4868 => x"3f",
          4869 => x"08",
          4870 => x"77",
          4871 => x"57",
          4872 => x"34",
          4873 => x"08",
          4874 => x"15",
          4875 => x"15",
          4876 => x"90",
          4877 => x"86",
          4878 => x"87",
          4879 => x"b6",
          4880 => x"b6",
          4881 => x"05",
          4882 => x"07",
          4883 => x"ff",
          4884 => x"2a",
          4885 => x"56",
          4886 => x"34",
          4887 => x"34",
          4888 => x"22",
          4889 => x"82",
          4890 => x"05",
          4891 => x"55",
          4892 => x"15",
          4893 => x"15",
          4894 => x"0d",
          4895 => x"0d",
          4896 => x"51",
          4897 => x"8f",
          4898 => x"83",
          4899 => x"70",
          4900 => x"06",
          4901 => x"70",
          4902 => x"0c",
          4903 => x"04",
          4904 => x"02",
          4905 => x"02",
          4906 => x"05",
          4907 => x"82",
          4908 => x"71",
          4909 => x"11",
          4910 => x"73",
          4911 => x"81",
          4912 => x"88",
          4913 => x"a4",
          4914 => x"22",
          4915 => x"ff",
          4916 => x"88",
          4917 => x"52",
          4918 => x"5b",
          4919 => x"55",
          4920 => x"70",
          4921 => x"82",
          4922 => x"14",
          4923 => x"52",
          4924 => x"15",
          4925 => x"15",
          4926 => x"90",
          4927 => x"70",
          4928 => x"33",
          4929 => x"07",
          4930 => x"8f",
          4931 => x"51",
          4932 => x"71",
          4933 => x"ff",
          4934 => x"88",
          4935 => x"51",
          4936 => x"34",
          4937 => x"06",
          4938 => x"12",
          4939 => x"90",
          4940 => x"71",
          4941 => x"81",
          4942 => x"3d",
          4943 => x"3d",
          4944 => x"90",
          4945 => x"05",
          4946 => x"70",
          4947 => x"11",
          4948 => x"87",
          4949 => x"8b",
          4950 => x"2b",
          4951 => x"59",
          4952 => x"72",
          4953 => x"33",
          4954 => x"71",
          4955 => x"70",
          4956 => x"56",
          4957 => x"84",
          4958 => x"85",
          4959 => x"b6",
          4960 => x"14",
          4961 => x"85",
          4962 => x"8b",
          4963 => x"2b",
          4964 => x"57",
          4965 => x"86",
          4966 => x"13",
          4967 => x"2b",
          4968 => x"2a",
          4969 => x"52",
          4970 => x"34",
          4971 => x"34",
          4972 => x"08",
          4973 => x"81",
          4974 => x"88",
          4975 => x"81",
          4976 => x"70",
          4977 => x"51",
          4978 => x"71",
          4979 => x"81",
          4980 => x"3d",
          4981 => x"3d",
          4982 => x"05",
          4983 => x"90",
          4984 => x"2b",
          4985 => x"33",
          4986 => x"71",
          4987 => x"70",
          4988 => x"70",
          4989 => x"33",
          4990 => x"71",
          4991 => x"53",
          4992 => x"52",
          4993 => x"53",
          4994 => x"25",
          4995 => x"72",
          4996 => x"3f",
          4997 => x"08",
          4998 => x"33",
          4999 => x"71",
          5000 => x"83",
          5001 => x"11",
          5002 => x"12",
          5003 => x"2b",
          5004 => x"2b",
          5005 => x"06",
          5006 => x"51",
          5007 => x"53",
          5008 => x"88",
          5009 => x"72",
          5010 => x"73",
          5011 => x"82",
          5012 => x"70",
          5013 => x"81",
          5014 => x"8b",
          5015 => x"2b",
          5016 => x"57",
          5017 => x"70",
          5018 => x"33",
          5019 => x"07",
          5020 => x"ff",
          5021 => x"2a",
          5022 => x"58",
          5023 => x"34",
          5024 => x"34",
          5025 => x"04",
          5026 => x"82",
          5027 => x"02",
          5028 => x"05",
          5029 => x"2b",
          5030 => x"11",
          5031 => x"33",
          5032 => x"71",
          5033 => x"59",
          5034 => x"56",
          5035 => x"71",
          5036 => x"33",
          5037 => x"07",
          5038 => x"a2",
          5039 => x"07",
          5040 => x"53",
          5041 => x"53",
          5042 => x"70",
          5043 => x"82",
          5044 => x"70",
          5045 => x"81",
          5046 => x"8b",
          5047 => x"2b",
          5048 => x"57",
          5049 => x"82",
          5050 => x"13",
          5051 => x"2b",
          5052 => x"2a",
          5053 => x"52",
          5054 => x"34",
          5055 => x"34",
          5056 => x"08",
          5057 => x"33",
          5058 => x"71",
          5059 => x"82",
          5060 => x"52",
          5061 => x"0d",
          5062 => x"0d",
          5063 => x"90",
          5064 => x"2a",
          5065 => x"ff",
          5066 => x"57",
          5067 => x"3f",
          5068 => x"08",
          5069 => x"71",
          5070 => x"33",
          5071 => x"71",
          5072 => x"83",
          5073 => x"11",
          5074 => x"12",
          5075 => x"2b",
          5076 => x"07",
          5077 => x"51",
          5078 => x"55",
          5079 => x"80",
          5080 => x"82",
          5081 => x"75",
          5082 => x"3f",
          5083 => x"84",
          5084 => x"15",
          5085 => x"2b",
          5086 => x"07",
          5087 => x"88",
          5088 => x"55",
          5089 => x"86",
          5090 => x"81",
          5091 => x"75",
          5092 => x"82",
          5093 => x"70",
          5094 => x"33",
          5095 => x"71",
          5096 => x"70",
          5097 => x"57",
          5098 => x"72",
          5099 => x"73",
          5100 => x"82",
          5101 => x"18",
          5102 => x"86",
          5103 => x"0b",
          5104 => x"82",
          5105 => x"53",
          5106 => x"34",
          5107 => x"34",
          5108 => x"08",
          5109 => x"81",
          5110 => x"88",
          5111 => x"82",
          5112 => x"70",
          5113 => x"51",
          5114 => x"74",
          5115 => x"81",
          5116 => x"3d",
          5117 => x"3d",
          5118 => x"82",
          5119 => x"84",
          5120 => x"3f",
          5121 => x"86",
          5122 => x"fe",
          5123 => x"3d",
          5124 => x"3d",
          5125 => x"52",
          5126 => x"3f",
          5127 => x"08",
          5128 => x"06",
          5129 => x"08",
          5130 => x"85",
          5131 => x"88",
          5132 => x"5f",
          5133 => x"5a",
          5134 => x"59",
          5135 => x"80",
          5136 => x"88",
          5137 => x"33",
          5138 => x"71",
          5139 => x"70",
          5140 => x"06",
          5141 => x"83",
          5142 => x"70",
          5143 => x"53",
          5144 => x"55",
          5145 => x"8a",
          5146 => x"2e",
          5147 => x"78",
          5148 => x"15",
          5149 => x"33",
          5150 => x"07",
          5151 => x"c2",
          5152 => x"ff",
          5153 => x"38",
          5154 => x"56",
          5155 => x"2b",
          5156 => x"08",
          5157 => x"81",
          5158 => x"88",
          5159 => x"81",
          5160 => x"51",
          5161 => x"5c",
          5162 => x"2e",
          5163 => x"55",
          5164 => x"78",
          5165 => x"38",
          5166 => x"80",
          5167 => x"38",
          5168 => x"09",
          5169 => x"38",
          5170 => x"f2",
          5171 => x"39",
          5172 => x"53",
          5173 => x"51",
          5174 => x"82",
          5175 => x"70",
          5176 => x"33",
          5177 => x"71",
          5178 => x"83",
          5179 => x"5a",
          5180 => x"05",
          5181 => x"83",
          5182 => x"70",
          5183 => x"59",
          5184 => x"84",
          5185 => x"81",
          5186 => x"76",
          5187 => x"82",
          5188 => x"75",
          5189 => x"11",
          5190 => x"11",
          5191 => x"33",
          5192 => x"07",
          5193 => x"53",
          5194 => x"5a",
          5195 => x"86",
          5196 => x"87",
          5197 => x"b6",
          5198 => x"1c",
          5199 => x"85",
          5200 => x"8b",
          5201 => x"2b",
          5202 => x"5a",
          5203 => x"54",
          5204 => x"34",
          5205 => x"34",
          5206 => x"08",
          5207 => x"1d",
          5208 => x"85",
          5209 => x"88",
          5210 => x"88",
          5211 => x"5f",
          5212 => x"73",
          5213 => x"75",
          5214 => x"82",
          5215 => x"1b",
          5216 => x"73",
          5217 => x"0c",
          5218 => x"04",
          5219 => x"74",
          5220 => x"90",
          5221 => x"f4",
          5222 => x"53",
          5223 => x"8b",
          5224 => x"fc",
          5225 => x"b6",
          5226 => x"72",
          5227 => x"0c",
          5228 => x"04",
          5229 => x"64",
          5230 => x"80",
          5231 => x"82",
          5232 => x"60",
          5233 => x"06",
          5234 => x"a9",
          5235 => x"38",
          5236 => x"b8",
          5237 => x"98",
          5238 => x"c7",
          5239 => x"38",
          5240 => x"92",
          5241 => x"83",
          5242 => x"51",
          5243 => x"82",
          5244 => x"83",
          5245 => x"82",
          5246 => x"7d",
          5247 => x"2a",
          5248 => x"ff",
          5249 => x"2b",
          5250 => x"33",
          5251 => x"71",
          5252 => x"70",
          5253 => x"83",
          5254 => x"70",
          5255 => x"05",
          5256 => x"1a",
          5257 => x"12",
          5258 => x"2b",
          5259 => x"2b",
          5260 => x"53",
          5261 => x"5c",
          5262 => x"5c",
          5263 => x"73",
          5264 => x"38",
          5265 => x"ff",
          5266 => x"70",
          5267 => x"06",
          5268 => x"16",
          5269 => x"33",
          5270 => x"07",
          5271 => x"1c",
          5272 => x"12",
          5273 => x"2b",
          5274 => x"07",
          5275 => x"52",
          5276 => x"80",
          5277 => x"78",
          5278 => x"83",
          5279 => x"41",
          5280 => x"27",
          5281 => x"60",
          5282 => x"7b",
          5283 => x"06",
          5284 => x"51",
          5285 => x"7a",
          5286 => x"06",
          5287 => x"39",
          5288 => x"7a",
          5289 => x"38",
          5290 => x"aa",
          5291 => x"39",
          5292 => x"7a",
          5293 => x"c8",
          5294 => x"82",
          5295 => x"12",
          5296 => x"2b",
          5297 => x"54",
          5298 => x"80",
          5299 => x"f7",
          5300 => x"b6",
          5301 => x"ff",
          5302 => x"54",
          5303 => x"83",
          5304 => x"90",
          5305 => x"05",
          5306 => x"ff",
          5307 => x"82",
          5308 => x"14",
          5309 => x"83",
          5310 => x"59",
          5311 => x"39",
          5312 => x"7a",
          5313 => x"d4",
          5314 => x"f5",
          5315 => x"b6",
          5316 => x"82",
          5317 => x"12",
          5318 => x"2b",
          5319 => x"54",
          5320 => x"80",
          5321 => x"f6",
          5322 => x"b6",
          5323 => x"ff",
          5324 => x"54",
          5325 => x"83",
          5326 => x"90",
          5327 => x"05",
          5328 => x"ff",
          5329 => x"82",
          5330 => x"14",
          5331 => x"62",
          5332 => x"5c",
          5333 => x"ff",
          5334 => x"39",
          5335 => x"54",
          5336 => x"82",
          5337 => x"5c",
          5338 => x"08",
          5339 => x"38",
          5340 => x"52",
          5341 => x"08",
          5342 => x"e9",
          5343 => x"f7",
          5344 => x"58",
          5345 => x"99",
          5346 => x"7a",
          5347 => x"f2",
          5348 => x"19",
          5349 => x"b6",
          5350 => x"84",
          5351 => x"f9",
          5352 => x"73",
          5353 => x"0c",
          5354 => x"04",
          5355 => x"77",
          5356 => x"52",
          5357 => x"3f",
          5358 => x"08",
          5359 => x"98",
          5360 => x"8e",
          5361 => x"80",
          5362 => x"98",
          5363 => x"9b",
          5364 => x"82",
          5365 => x"86",
          5366 => x"ff",
          5367 => x"8f",
          5368 => x"81",
          5369 => x"26",
          5370 => x"b6",
          5371 => x"52",
          5372 => x"98",
          5373 => x"0d",
          5374 => x"0d",
          5375 => x"33",
          5376 => x"9f",
          5377 => x"53",
          5378 => x"81",
          5379 => x"38",
          5380 => x"87",
          5381 => x"11",
          5382 => x"54",
          5383 => x"84",
          5384 => x"54",
          5385 => x"87",
          5386 => x"11",
          5387 => x"0c",
          5388 => x"c0",
          5389 => x"70",
          5390 => x"70",
          5391 => x"51",
          5392 => x"8a",
          5393 => x"98",
          5394 => x"70",
          5395 => x"08",
          5396 => x"06",
          5397 => x"38",
          5398 => x"8c",
          5399 => x"80",
          5400 => x"71",
          5401 => x"14",
          5402 => x"94",
          5403 => x"70",
          5404 => x"0c",
          5405 => x"04",
          5406 => x"60",
          5407 => x"8c",
          5408 => x"33",
          5409 => x"5b",
          5410 => x"5a",
          5411 => x"82",
          5412 => x"81",
          5413 => x"52",
          5414 => x"38",
          5415 => x"84",
          5416 => x"92",
          5417 => x"c0",
          5418 => x"87",
          5419 => x"13",
          5420 => x"57",
          5421 => x"0b",
          5422 => x"8c",
          5423 => x"0c",
          5424 => x"75",
          5425 => x"2a",
          5426 => x"51",
          5427 => x"80",
          5428 => x"7b",
          5429 => x"7b",
          5430 => x"5d",
          5431 => x"59",
          5432 => x"06",
          5433 => x"73",
          5434 => x"81",
          5435 => x"ff",
          5436 => x"72",
          5437 => x"38",
          5438 => x"8c",
          5439 => x"c3",
          5440 => x"98",
          5441 => x"71",
          5442 => x"38",
          5443 => x"2e",
          5444 => x"76",
          5445 => x"92",
          5446 => x"72",
          5447 => x"06",
          5448 => x"f7",
          5449 => x"5a",
          5450 => x"80",
          5451 => x"70",
          5452 => x"5a",
          5453 => x"80",
          5454 => x"73",
          5455 => x"06",
          5456 => x"38",
          5457 => x"fe",
          5458 => x"fc",
          5459 => x"52",
          5460 => x"83",
          5461 => x"71",
          5462 => x"b6",
          5463 => x"3d",
          5464 => x"3d",
          5465 => x"64",
          5466 => x"bf",
          5467 => x"40",
          5468 => x"59",
          5469 => x"58",
          5470 => x"82",
          5471 => x"81",
          5472 => x"52",
          5473 => x"09",
          5474 => x"b1",
          5475 => x"84",
          5476 => x"92",
          5477 => x"c0",
          5478 => x"87",
          5479 => x"13",
          5480 => x"56",
          5481 => x"87",
          5482 => x"0c",
          5483 => x"82",
          5484 => x"58",
          5485 => x"84",
          5486 => x"06",
          5487 => x"71",
          5488 => x"38",
          5489 => x"05",
          5490 => x"0c",
          5491 => x"73",
          5492 => x"81",
          5493 => x"71",
          5494 => x"38",
          5495 => x"8c",
          5496 => x"d0",
          5497 => x"98",
          5498 => x"71",
          5499 => x"38",
          5500 => x"2e",
          5501 => x"76",
          5502 => x"92",
          5503 => x"72",
          5504 => x"06",
          5505 => x"f7",
          5506 => x"59",
          5507 => x"1a",
          5508 => x"06",
          5509 => x"59",
          5510 => x"80",
          5511 => x"73",
          5512 => x"06",
          5513 => x"38",
          5514 => x"fe",
          5515 => x"fc",
          5516 => x"52",
          5517 => x"83",
          5518 => x"71",
          5519 => x"b6",
          5520 => x"3d",
          5521 => x"3d",
          5522 => x"84",
          5523 => x"33",
          5524 => x"a7",
          5525 => x"54",
          5526 => x"fa",
          5527 => x"b6",
          5528 => x"06",
          5529 => x"72",
          5530 => x"85",
          5531 => x"98",
          5532 => x"56",
          5533 => x"80",
          5534 => x"76",
          5535 => x"74",
          5536 => x"c0",
          5537 => x"54",
          5538 => x"2e",
          5539 => x"d4",
          5540 => x"2e",
          5541 => x"80",
          5542 => x"08",
          5543 => x"70",
          5544 => x"51",
          5545 => x"2e",
          5546 => x"c0",
          5547 => x"52",
          5548 => x"87",
          5549 => x"08",
          5550 => x"38",
          5551 => x"87",
          5552 => x"14",
          5553 => x"70",
          5554 => x"52",
          5555 => x"96",
          5556 => x"92",
          5557 => x"0a",
          5558 => x"39",
          5559 => x"0c",
          5560 => x"39",
          5561 => x"54",
          5562 => x"98",
          5563 => x"0d",
          5564 => x"0d",
          5565 => x"33",
          5566 => x"88",
          5567 => x"b6",
          5568 => x"51",
          5569 => x"04",
          5570 => x"75",
          5571 => x"82",
          5572 => x"90",
          5573 => x"2b",
          5574 => x"33",
          5575 => x"88",
          5576 => x"71",
          5577 => x"98",
          5578 => x"54",
          5579 => x"85",
          5580 => x"ff",
          5581 => x"02",
          5582 => x"05",
          5583 => x"70",
          5584 => x"05",
          5585 => x"88",
          5586 => x"72",
          5587 => x"0d",
          5588 => x"0d",
          5589 => x"52",
          5590 => x"81",
          5591 => x"70",
          5592 => x"70",
          5593 => x"05",
          5594 => x"88",
          5595 => x"72",
          5596 => x"54",
          5597 => x"2a",
          5598 => x"34",
          5599 => x"04",
          5600 => x"76",
          5601 => x"54",
          5602 => x"2e",
          5603 => x"70",
          5604 => x"33",
          5605 => x"05",
          5606 => x"11",
          5607 => x"84",
          5608 => x"fe",
          5609 => x"77",
          5610 => x"53",
          5611 => x"81",
          5612 => x"ff",
          5613 => x"f4",
          5614 => x"0d",
          5615 => x"0d",
          5616 => x"56",
          5617 => x"70",
          5618 => x"33",
          5619 => x"05",
          5620 => x"71",
          5621 => x"56",
          5622 => x"72",
          5623 => x"38",
          5624 => x"e2",
          5625 => x"b6",
          5626 => x"3d",
          5627 => x"3d",
          5628 => x"54",
          5629 => x"71",
          5630 => x"38",
          5631 => x"70",
          5632 => x"f3",
          5633 => x"82",
          5634 => x"84",
          5635 => x"80",
          5636 => x"98",
          5637 => x"0b",
          5638 => x"0c",
          5639 => x"0d",
          5640 => x"0b",
          5641 => x"56",
          5642 => x"2e",
          5643 => x"81",
          5644 => x"08",
          5645 => x"70",
          5646 => x"33",
          5647 => x"a2",
          5648 => x"98",
          5649 => x"09",
          5650 => x"38",
          5651 => x"08",
          5652 => x"b0",
          5653 => x"a4",
          5654 => x"9c",
          5655 => x"56",
          5656 => x"27",
          5657 => x"16",
          5658 => x"82",
          5659 => x"06",
          5660 => x"54",
          5661 => x"78",
          5662 => x"33",
          5663 => x"3f",
          5664 => x"5a",
          5665 => x"98",
          5666 => x"0d",
          5667 => x"0d",
          5668 => x"56",
          5669 => x"b0",
          5670 => x"af",
          5671 => x"fe",
          5672 => x"b6",
          5673 => x"82",
          5674 => x"9f",
          5675 => x"74",
          5676 => x"52",
          5677 => x"51",
          5678 => x"82",
          5679 => x"80",
          5680 => x"ff",
          5681 => x"74",
          5682 => x"76",
          5683 => x"0c",
          5684 => x"04",
          5685 => x"7a",
          5686 => x"fe",
          5687 => x"b6",
          5688 => x"82",
          5689 => x"81",
          5690 => x"33",
          5691 => x"2e",
          5692 => x"80",
          5693 => x"17",
          5694 => x"81",
          5695 => x"06",
          5696 => x"84",
          5697 => x"b6",
          5698 => x"b4",
          5699 => x"56",
          5700 => x"82",
          5701 => x"84",
          5702 => x"fc",
          5703 => x"8b",
          5704 => x"52",
          5705 => x"a9",
          5706 => x"85",
          5707 => x"84",
          5708 => x"fc",
          5709 => x"17",
          5710 => x"9c",
          5711 => x"91",
          5712 => x"08",
          5713 => x"17",
          5714 => x"3f",
          5715 => x"81",
          5716 => x"19",
          5717 => x"53",
          5718 => x"17",
          5719 => x"82",
          5720 => x"18",
          5721 => x"80",
          5722 => x"33",
          5723 => x"3f",
          5724 => x"08",
          5725 => x"38",
          5726 => x"82",
          5727 => x"8a",
          5728 => x"fb",
          5729 => x"fe",
          5730 => x"08",
          5731 => x"56",
          5732 => x"74",
          5733 => x"38",
          5734 => x"75",
          5735 => x"16",
          5736 => x"53",
          5737 => x"98",
          5738 => x"0d",
          5739 => x"0d",
          5740 => x"08",
          5741 => x"81",
          5742 => x"df",
          5743 => x"15",
          5744 => x"d7",
          5745 => x"33",
          5746 => x"82",
          5747 => x"38",
          5748 => x"89",
          5749 => x"2e",
          5750 => x"bf",
          5751 => x"2e",
          5752 => x"81",
          5753 => x"81",
          5754 => x"89",
          5755 => x"08",
          5756 => x"52",
          5757 => x"3f",
          5758 => x"08",
          5759 => x"74",
          5760 => x"14",
          5761 => x"81",
          5762 => x"2a",
          5763 => x"05",
          5764 => x"57",
          5765 => x"f5",
          5766 => x"98",
          5767 => x"38",
          5768 => x"06",
          5769 => x"33",
          5770 => x"78",
          5771 => x"06",
          5772 => x"5c",
          5773 => x"53",
          5774 => x"38",
          5775 => x"06",
          5776 => x"39",
          5777 => x"a4",
          5778 => x"52",
          5779 => x"bd",
          5780 => x"98",
          5781 => x"38",
          5782 => x"fe",
          5783 => x"b4",
          5784 => x"8d",
          5785 => x"98",
          5786 => x"ff",
          5787 => x"39",
          5788 => x"a4",
          5789 => x"52",
          5790 => x"91",
          5791 => x"98",
          5792 => x"76",
          5793 => x"fc",
          5794 => x"b4",
          5795 => x"f8",
          5796 => x"98",
          5797 => x"06",
          5798 => x"81",
          5799 => x"b6",
          5800 => x"3d",
          5801 => x"3d",
          5802 => x"7e",
          5803 => x"82",
          5804 => x"27",
          5805 => x"76",
          5806 => x"27",
          5807 => x"75",
          5808 => x"79",
          5809 => x"38",
          5810 => x"89",
          5811 => x"2e",
          5812 => x"80",
          5813 => x"2e",
          5814 => x"81",
          5815 => x"81",
          5816 => x"89",
          5817 => x"08",
          5818 => x"52",
          5819 => x"3f",
          5820 => x"08",
          5821 => x"98",
          5822 => x"38",
          5823 => x"06",
          5824 => x"81",
          5825 => x"06",
          5826 => x"77",
          5827 => x"2e",
          5828 => x"84",
          5829 => x"06",
          5830 => x"06",
          5831 => x"53",
          5832 => x"81",
          5833 => x"34",
          5834 => x"a4",
          5835 => x"52",
          5836 => x"d9",
          5837 => x"98",
          5838 => x"b6",
          5839 => x"94",
          5840 => x"ff",
          5841 => x"05",
          5842 => x"54",
          5843 => x"38",
          5844 => x"74",
          5845 => x"06",
          5846 => x"07",
          5847 => x"74",
          5848 => x"39",
          5849 => x"a4",
          5850 => x"52",
          5851 => x"9d",
          5852 => x"98",
          5853 => x"b6",
          5854 => x"d8",
          5855 => x"ff",
          5856 => x"76",
          5857 => x"06",
          5858 => x"05",
          5859 => x"3f",
          5860 => x"87",
          5861 => x"08",
          5862 => x"51",
          5863 => x"82",
          5864 => x"59",
          5865 => x"08",
          5866 => x"f0",
          5867 => x"82",
          5868 => x"06",
          5869 => x"05",
          5870 => x"54",
          5871 => x"3f",
          5872 => x"08",
          5873 => x"74",
          5874 => x"51",
          5875 => x"81",
          5876 => x"34",
          5877 => x"98",
          5878 => x"0d",
          5879 => x"0d",
          5880 => x"72",
          5881 => x"56",
          5882 => x"27",
          5883 => x"98",
          5884 => x"9d",
          5885 => x"2e",
          5886 => x"53",
          5887 => x"51",
          5888 => x"82",
          5889 => x"54",
          5890 => x"08",
          5891 => x"93",
          5892 => x"80",
          5893 => x"54",
          5894 => x"82",
          5895 => x"54",
          5896 => x"74",
          5897 => x"fb",
          5898 => x"b6",
          5899 => x"82",
          5900 => x"80",
          5901 => x"38",
          5902 => x"08",
          5903 => x"38",
          5904 => x"08",
          5905 => x"38",
          5906 => x"52",
          5907 => x"d6",
          5908 => x"98",
          5909 => x"98",
          5910 => x"11",
          5911 => x"57",
          5912 => x"74",
          5913 => x"81",
          5914 => x"0c",
          5915 => x"81",
          5916 => x"84",
          5917 => x"55",
          5918 => x"ff",
          5919 => x"54",
          5920 => x"98",
          5921 => x"0d",
          5922 => x"0d",
          5923 => x"08",
          5924 => x"79",
          5925 => x"17",
          5926 => x"80",
          5927 => x"98",
          5928 => x"26",
          5929 => x"58",
          5930 => x"52",
          5931 => x"fd",
          5932 => x"74",
          5933 => x"08",
          5934 => x"38",
          5935 => x"08",
          5936 => x"98",
          5937 => x"82",
          5938 => x"17",
          5939 => x"98",
          5940 => x"c7",
          5941 => x"90",
          5942 => x"56",
          5943 => x"2e",
          5944 => x"77",
          5945 => x"81",
          5946 => x"38",
          5947 => x"98",
          5948 => x"26",
          5949 => x"56",
          5950 => x"51",
          5951 => x"80",
          5952 => x"98",
          5953 => x"09",
          5954 => x"38",
          5955 => x"08",
          5956 => x"98",
          5957 => x"30",
          5958 => x"80",
          5959 => x"07",
          5960 => x"08",
          5961 => x"55",
          5962 => x"ef",
          5963 => x"98",
          5964 => x"95",
          5965 => x"08",
          5966 => x"27",
          5967 => x"98",
          5968 => x"89",
          5969 => x"85",
          5970 => x"db",
          5971 => x"81",
          5972 => x"17",
          5973 => x"89",
          5974 => x"75",
          5975 => x"ac",
          5976 => x"7a",
          5977 => x"3f",
          5978 => x"08",
          5979 => x"38",
          5980 => x"b6",
          5981 => x"2e",
          5982 => x"86",
          5983 => x"98",
          5984 => x"b6",
          5985 => x"70",
          5986 => x"07",
          5987 => x"7c",
          5988 => x"55",
          5989 => x"f8",
          5990 => x"2e",
          5991 => x"ff",
          5992 => x"55",
          5993 => x"ff",
          5994 => x"76",
          5995 => x"3f",
          5996 => x"08",
          5997 => x"08",
          5998 => x"b6",
          5999 => x"80",
          6000 => x"55",
          6001 => x"94",
          6002 => x"2e",
          6003 => x"53",
          6004 => x"51",
          6005 => x"82",
          6006 => x"55",
          6007 => x"75",
          6008 => x"98",
          6009 => x"05",
          6010 => x"56",
          6011 => x"26",
          6012 => x"15",
          6013 => x"84",
          6014 => x"07",
          6015 => x"18",
          6016 => x"ff",
          6017 => x"2e",
          6018 => x"39",
          6019 => x"39",
          6020 => x"08",
          6021 => x"81",
          6022 => x"74",
          6023 => x"0c",
          6024 => x"04",
          6025 => x"7a",
          6026 => x"f3",
          6027 => x"b6",
          6028 => x"81",
          6029 => x"98",
          6030 => x"38",
          6031 => x"51",
          6032 => x"82",
          6033 => x"82",
          6034 => x"b0",
          6035 => x"84",
          6036 => x"52",
          6037 => x"52",
          6038 => x"3f",
          6039 => x"39",
          6040 => x"8a",
          6041 => x"75",
          6042 => x"38",
          6043 => x"19",
          6044 => x"81",
          6045 => x"ed",
          6046 => x"b6",
          6047 => x"2e",
          6048 => x"15",
          6049 => x"70",
          6050 => x"07",
          6051 => x"53",
          6052 => x"75",
          6053 => x"0c",
          6054 => x"04",
          6055 => x"7a",
          6056 => x"58",
          6057 => x"f0",
          6058 => x"80",
          6059 => x"9f",
          6060 => x"80",
          6061 => x"90",
          6062 => x"17",
          6063 => x"aa",
          6064 => x"53",
          6065 => x"88",
          6066 => x"08",
          6067 => x"38",
          6068 => x"53",
          6069 => x"17",
          6070 => x"72",
          6071 => x"fe",
          6072 => x"08",
          6073 => x"80",
          6074 => x"16",
          6075 => x"2b",
          6076 => x"75",
          6077 => x"73",
          6078 => x"f5",
          6079 => x"b6",
          6080 => x"82",
          6081 => x"ff",
          6082 => x"81",
          6083 => x"98",
          6084 => x"38",
          6085 => x"82",
          6086 => x"26",
          6087 => x"58",
          6088 => x"73",
          6089 => x"39",
          6090 => x"51",
          6091 => x"82",
          6092 => x"98",
          6093 => x"94",
          6094 => x"17",
          6095 => x"58",
          6096 => x"9a",
          6097 => x"81",
          6098 => x"74",
          6099 => x"98",
          6100 => x"83",
          6101 => x"b4",
          6102 => x"0c",
          6103 => x"82",
          6104 => x"8a",
          6105 => x"f8",
          6106 => x"70",
          6107 => x"08",
          6108 => x"57",
          6109 => x"0a",
          6110 => x"38",
          6111 => x"15",
          6112 => x"08",
          6113 => x"72",
          6114 => x"cb",
          6115 => x"ff",
          6116 => x"81",
          6117 => x"13",
          6118 => x"94",
          6119 => x"74",
          6120 => x"85",
          6121 => x"22",
          6122 => x"73",
          6123 => x"38",
          6124 => x"8a",
          6125 => x"05",
          6126 => x"06",
          6127 => x"8a",
          6128 => x"73",
          6129 => x"3f",
          6130 => x"08",
          6131 => x"81",
          6132 => x"98",
          6133 => x"ff",
          6134 => x"82",
          6135 => x"ff",
          6136 => x"38",
          6137 => x"82",
          6138 => x"26",
          6139 => x"7b",
          6140 => x"98",
          6141 => x"55",
          6142 => x"94",
          6143 => x"73",
          6144 => x"3f",
          6145 => x"08",
          6146 => x"82",
          6147 => x"80",
          6148 => x"38",
          6149 => x"b6",
          6150 => x"2e",
          6151 => x"55",
          6152 => x"08",
          6153 => x"38",
          6154 => x"08",
          6155 => x"fb",
          6156 => x"b6",
          6157 => x"38",
          6158 => x"0c",
          6159 => x"51",
          6160 => x"82",
          6161 => x"98",
          6162 => x"90",
          6163 => x"16",
          6164 => x"15",
          6165 => x"74",
          6166 => x"0c",
          6167 => x"04",
          6168 => x"7b",
          6169 => x"5b",
          6170 => x"52",
          6171 => x"ac",
          6172 => x"98",
          6173 => x"b6",
          6174 => x"ec",
          6175 => x"98",
          6176 => x"17",
          6177 => x"51",
          6178 => x"82",
          6179 => x"54",
          6180 => x"08",
          6181 => x"82",
          6182 => x"9c",
          6183 => x"33",
          6184 => x"72",
          6185 => x"09",
          6186 => x"38",
          6187 => x"b6",
          6188 => x"72",
          6189 => x"55",
          6190 => x"53",
          6191 => x"8e",
          6192 => x"56",
          6193 => x"09",
          6194 => x"38",
          6195 => x"b6",
          6196 => x"81",
          6197 => x"fd",
          6198 => x"b6",
          6199 => x"82",
          6200 => x"80",
          6201 => x"38",
          6202 => x"09",
          6203 => x"38",
          6204 => x"82",
          6205 => x"8b",
          6206 => x"fd",
          6207 => x"9a",
          6208 => x"eb",
          6209 => x"b6",
          6210 => x"ff",
          6211 => x"70",
          6212 => x"53",
          6213 => x"09",
          6214 => x"38",
          6215 => x"eb",
          6216 => x"b6",
          6217 => x"2b",
          6218 => x"72",
          6219 => x"0c",
          6220 => x"04",
          6221 => x"77",
          6222 => x"ff",
          6223 => x"9a",
          6224 => x"55",
          6225 => x"76",
          6226 => x"53",
          6227 => x"09",
          6228 => x"38",
          6229 => x"52",
          6230 => x"eb",
          6231 => x"3d",
          6232 => x"3d",
          6233 => x"5b",
          6234 => x"08",
          6235 => x"15",
          6236 => x"81",
          6237 => x"15",
          6238 => x"51",
          6239 => x"82",
          6240 => x"58",
          6241 => x"08",
          6242 => x"9c",
          6243 => x"33",
          6244 => x"86",
          6245 => x"80",
          6246 => x"13",
          6247 => x"06",
          6248 => x"06",
          6249 => x"72",
          6250 => x"82",
          6251 => x"53",
          6252 => x"2e",
          6253 => x"53",
          6254 => x"a9",
          6255 => x"74",
          6256 => x"72",
          6257 => x"38",
          6258 => x"99",
          6259 => x"98",
          6260 => x"06",
          6261 => x"88",
          6262 => x"06",
          6263 => x"54",
          6264 => x"a0",
          6265 => x"74",
          6266 => x"3f",
          6267 => x"08",
          6268 => x"98",
          6269 => x"98",
          6270 => x"fa",
          6271 => x"80",
          6272 => x"0c",
          6273 => x"98",
          6274 => x"0d",
          6275 => x"0d",
          6276 => x"57",
          6277 => x"73",
          6278 => x"3f",
          6279 => x"08",
          6280 => x"98",
          6281 => x"98",
          6282 => x"75",
          6283 => x"3f",
          6284 => x"08",
          6285 => x"98",
          6286 => x"a0",
          6287 => x"98",
          6288 => x"14",
          6289 => x"db",
          6290 => x"a0",
          6291 => x"14",
          6292 => x"ac",
          6293 => x"83",
          6294 => x"82",
          6295 => x"87",
          6296 => x"fd",
          6297 => x"70",
          6298 => x"08",
          6299 => x"55",
          6300 => x"3f",
          6301 => x"08",
          6302 => x"13",
          6303 => x"73",
          6304 => x"83",
          6305 => x"3d",
          6306 => x"3d",
          6307 => x"57",
          6308 => x"89",
          6309 => x"17",
          6310 => x"81",
          6311 => x"70",
          6312 => x"55",
          6313 => x"08",
          6314 => x"81",
          6315 => x"52",
          6316 => x"a8",
          6317 => x"2e",
          6318 => x"84",
          6319 => x"52",
          6320 => x"09",
          6321 => x"38",
          6322 => x"81",
          6323 => x"81",
          6324 => x"73",
          6325 => x"55",
          6326 => x"55",
          6327 => x"c5",
          6328 => x"88",
          6329 => x"0b",
          6330 => x"9c",
          6331 => x"8b",
          6332 => x"17",
          6333 => x"08",
          6334 => x"52",
          6335 => x"82",
          6336 => x"76",
          6337 => x"51",
          6338 => x"82",
          6339 => x"86",
          6340 => x"12",
          6341 => x"3f",
          6342 => x"08",
          6343 => x"88",
          6344 => x"f3",
          6345 => x"70",
          6346 => x"80",
          6347 => x"51",
          6348 => x"af",
          6349 => x"81",
          6350 => x"dc",
          6351 => x"74",
          6352 => x"38",
          6353 => x"88",
          6354 => x"39",
          6355 => x"80",
          6356 => x"56",
          6357 => x"af",
          6358 => x"06",
          6359 => x"56",
          6360 => x"32",
          6361 => x"80",
          6362 => x"51",
          6363 => x"dc",
          6364 => x"1c",
          6365 => x"33",
          6366 => x"9f",
          6367 => x"ff",
          6368 => x"1c",
          6369 => x"7a",
          6370 => x"3f",
          6371 => x"08",
          6372 => x"39",
          6373 => x"a0",
          6374 => x"5e",
          6375 => x"52",
          6376 => x"ff",
          6377 => x"59",
          6378 => x"33",
          6379 => x"ae",
          6380 => x"06",
          6381 => x"78",
          6382 => x"81",
          6383 => x"32",
          6384 => x"9f",
          6385 => x"26",
          6386 => x"53",
          6387 => x"73",
          6388 => x"17",
          6389 => x"34",
          6390 => x"db",
          6391 => x"32",
          6392 => x"9f",
          6393 => x"54",
          6394 => x"2e",
          6395 => x"80",
          6396 => x"75",
          6397 => x"bd",
          6398 => x"7e",
          6399 => x"a0",
          6400 => x"bd",
          6401 => x"82",
          6402 => x"18",
          6403 => x"1a",
          6404 => x"a0",
          6405 => x"fc",
          6406 => x"32",
          6407 => x"80",
          6408 => x"30",
          6409 => x"71",
          6410 => x"51",
          6411 => x"55",
          6412 => x"ac",
          6413 => x"81",
          6414 => x"78",
          6415 => x"51",
          6416 => x"af",
          6417 => x"06",
          6418 => x"55",
          6419 => x"32",
          6420 => x"80",
          6421 => x"51",
          6422 => x"db",
          6423 => x"39",
          6424 => x"09",
          6425 => x"38",
          6426 => x"7c",
          6427 => x"54",
          6428 => x"a2",
          6429 => x"32",
          6430 => x"ae",
          6431 => x"72",
          6432 => x"9f",
          6433 => x"51",
          6434 => x"74",
          6435 => x"88",
          6436 => x"fe",
          6437 => x"98",
          6438 => x"80",
          6439 => x"75",
          6440 => x"82",
          6441 => x"33",
          6442 => x"51",
          6443 => x"82",
          6444 => x"80",
          6445 => x"78",
          6446 => x"81",
          6447 => x"5a",
          6448 => x"d2",
          6449 => x"98",
          6450 => x"80",
          6451 => x"1c",
          6452 => x"27",
          6453 => x"79",
          6454 => x"74",
          6455 => x"7a",
          6456 => x"74",
          6457 => x"39",
          6458 => x"af",
          6459 => x"fe",
          6460 => x"98",
          6461 => x"ff",
          6462 => x"73",
          6463 => x"38",
          6464 => x"81",
          6465 => x"54",
          6466 => x"75",
          6467 => x"17",
          6468 => x"39",
          6469 => x"0c",
          6470 => x"99",
          6471 => x"54",
          6472 => x"2e",
          6473 => x"84",
          6474 => x"34",
          6475 => x"76",
          6476 => x"8b",
          6477 => x"81",
          6478 => x"56",
          6479 => x"80",
          6480 => x"1b",
          6481 => x"08",
          6482 => x"51",
          6483 => x"82",
          6484 => x"56",
          6485 => x"08",
          6486 => x"98",
          6487 => x"76",
          6488 => x"3f",
          6489 => x"08",
          6490 => x"98",
          6491 => x"38",
          6492 => x"70",
          6493 => x"73",
          6494 => x"be",
          6495 => x"33",
          6496 => x"73",
          6497 => x"8b",
          6498 => x"83",
          6499 => x"06",
          6500 => x"73",
          6501 => x"53",
          6502 => x"51",
          6503 => x"82",
          6504 => x"80",
          6505 => x"75",
          6506 => x"f3",
          6507 => x"9f",
          6508 => x"1c",
          6509 => x"74",
          6510 => x"38",
          6511 => x"09",
          6512 => x"e7",
          6513 => x"2a",
          6514 => x"77",
          6515 => x"51",
          6516 => x"2e",
          6517 => x"81",
          6518 => x"80",
          6519 => x"38",
          6520 => x"ab",
          6521 => x"55",
          6522 => x"75",
          6523 => x"73",
          6524 => x"55",
          6525 => x"82",
          6526 => x"06",
          6527 => x"ab",
          6528 => x"33",
          6529 => x"70",
          6530 => x"55",
          6531 => x"2e",
          6532 => x"1b",
          6533 => x"06",
          6534 => x"52",
          6535 => x"db",
          6536 => x"98",
          6537 => x"0c",
          6538 => x"74",
          6539 => x"0c",
          6540 => x"04",
          6541 => x"7c",
          6542 => x"08",
          6543 => x"55",
          6544 => x"59",
          6545 => x"81",
          6546 => x"70",
          6547 => x"33",
          6548 => x"52",
          6549 => x"2e",
          6550 => x"ee",
          6551 => x"2e",
          6552 => x"81",
          6553 => x"33",
          6554 => x"81",
          6555 => x"52",
          6556 => x"26",
          6557 => x"14",
          6558 => x"06",
          6559 => x"52",
          6560 => x"80",
          6561 => x"0b",
          6562 => x"59",
          6563 => x"7a",
          6564 => x"70",
          6565 => x"33",
          6566 => x"05",
          6567 => x"9f",
          6568 => x"53",
          6569 => x"89",
          6570 => x"70",
          6571 => x"54",
          6572 => x"12",
          6573 => x"26",
          6574 => x"12",
          6575 => x"06",
          6576 => x"30",
          6577 => x"51",
          6578 => x"2e",
          6579 => x"85",
          6580 => x"be",
          6581 => x"74",
          6582 => x"30",
          6583 => x"9f",
          6584 => x"2a",
          6585 => x"54",
          6586 => x"2e",
          6587 => x"15",
          6588 => x"55",
          6589 => x"ff",
          6590 => x"39",
          6591 => x"86",
          6592 => x"7c",
          6593 => x"51",
          6594 => x"cd",
          6595 => x"70",
          6596 => x"0c",
          6597 => x"04",
          6598 => x"78",
          6599 => x"83",
          6600 => x"0b",
          6601 => x"79",
          6602 => x"e2",
          6603 => x"55",
          6604 => x"08",
          6605 => x"84",
          6606 => x"df",
          6607 => x"b6",
          6608 => x"ff",
          6609 => x"83",
          6610 => x"d4",
          6611 => x"81",
          6612 => x"38",
          6613 => x"17",
          6614 => x"74",
          6615 => x"09",
          6616 => x"38",
          6617 => x"81",
          6618 => x"30",
          6619 => x"79",
          6620 => x"54",
          6621 => x"74",
          6622 => x"09",
          6623 => x"38",
          6624 => x"af",
          6625 => x"ea",
          6626 => x"b1",
          6627 => x"98",
          6628 => x"b6",
          6629 => x"2e",
          6630 => x"53",
          6631 => x"52",
          6632 => x"51",
          6633 => x"82",
          6634 => x"55",
          6635 => x"08",
          6636 => x"38",
          6637 => x"82",
          6638 => x"88",
          6639 => x"f2",
          6640 => x"02",
          6641 => x"cb",
          6642 => x"55",
          6643 => x"60",
          6644 => x"3f",
          6645 => x"08",
          6646 => x"80",
          6647 => x"98",
          6648 => x"fc",
          6649 => x"98",
          6650 => x"82",
          6651 => x"70",
          6652 => x"8c",
          6653 => x"2e",
          6654 => x"73",
          6655 => x"81",
          6656 => x"33",
          6657 => x"80",
          6658 => x"81",
          6659 => x"d7",
          6660 => x"b6",
          6661 => x"ff",
          6662 => x"06",
          6663 => x"98",
          6664 => x"2e",
          6665 => x"74",
          6666 => x"81",
          6667 => x"8a",
          6668 => x"ac",
          6669 => x"39",
          6670 => x"77",
          6671 => x"81",
          6672 => x"33",
          6673 => x"3f",
          6674 => x"08",
          6675 => x"70",
          6676 => x"55",
          6677 => x"86",
          6678 => x"80",
          6679 => x"74",
          6680 => x"81",
          6681 => x"8a",
          6682 => x"f4",
          6683 => x"53",
          6684 => x"fd",
          6685 => x"b6",
          6686 => x"ff",
          6687 => x"82",
          6688 => x"06",
          6689 => x"8c",
          6690 => x"58",
          6691 => x"f6",
          6692 => x"58",
          6693 => x"2e",
          6694 => x"fa",
          6695 => x"e8",
          6696 => x"98",
          6697 => x"78",
          6698 => x"5a",
          6699 => x"90",
          6700 => x"75",
          6701 => x"38",
          6702 => x"3d",
          6703 => x"70",
          6704 => x"08",
          6705 => x"7a",
          6706 => x"38",
          6707 => x"51",
          6708 => x"82",
          6709 => x"81",
          6710 => x"81",
          6711 => x"38",
          6712 => x"83",
          6713 => x"38",
          6714 => x"84",
          6715 => x"38",
          6716 => x"81",
          6717 => x"38",
          6718 => x"db",
          6719 => x"b6",
          6720 => x"ff",
          6721 => x"72",
          6722 => x"09",
          6723 => x"d0",
          6724 => x"14",
          6725 => x"3f",
          6726 => x"08",
          6727 => x"06",
          6728 => x"38",
          6729 => x"51",
          6730 => x"82",
          6731 => x"58",
          6732 => x"0c",
          6733 => x"33",
          6734 => x"80",
          6735 => x"ff",
          6736 => x"ff",
          6737 => x"55",
          6738 => x"81",
          6739 => x"38",
          6740 => x"06",
          6741 => x"80",
          6742 => x"52",
          6743 => x"8a",
          6744 => x"80",
          6745 => x"ff",
          6746 => x"53",
          6747 => x"86",
          6748 => x"83",
          6749 => x"c5",
          6750 => x"f5",
          6751 => x"98",
          6752 => x"b6",
          6753 => x"15",
          6754 => x"06",
          6755 => x"76",
          6756 => x"80",
          6757 => x"da",
          6758 => x"b6",
          6759 => x"ff",
          6760 => x"74",
          6761 => x"d4",
          6762 => x"dc",
          6763 => x"98",
          6764 => x"c2",
          6765 => x"b9",
          6766 => x"98",
          6767 => x"ff",
          6768 => x"56",
          6769 => x"83",
          6770 => x"14",
          6771 => x"71",
          6772 => x"5a",
          6773 => x"26",
          6774 => x"8a",
          6775 => x"74",
          6776 => x"fe",
          6777 => x"82",
          6778 => x"55",
          6779 => x"08",
          6780 => x"ec",
          6781 => x"98",
          6782 => x"ff",
          6783 => x"83",
          6784 => x"74",
          6785 => x"26",
          6786 => x"57",
          6787 => x"26",
          6788 => x"57",
          6789 => x"56",
          6790 => x"82",
          6791 => x"15",
          6792 => x"0c",
          6793 => x"0c",
          6794 => x"a4",
          6795 => x"1d",
          6796 => x"54",
          6797 => x"2e",
          6798 => x"af",
          6799 => x"14",
          6800 => x"3f",
          6801 => x"08",
          6802 => x"06",
          6803 => x"72",
          6804 => x"79",
          6805 => x"80",
          6806 => x"d9",
          6807 => x"b6",
          6808 => x"15",
          6809 => x"2b",
          6810 => x"8d",
          6811 => x"2e",
          6812 => x"77",
          6813 => x"0c",
          6814 => x"76",
          6815 => x"38",
          6816 => x"70",
          6817 => x"81",
          6818 => x"53",
          6819 => x"89",
          6820 => x"56",
          6821 => x"08",
          6822 => x"38",
          6823 => x"15",
          6824 => x"8c",
          6825 => x"80",
          6826 => x"34",
          6827 => x"09",
          6828 => x"92",
          6829 => x"14",
          6830 => x"3f",
          6831 => x"08",
          6832 => x"06",
          6833 => x"2e",
          6834 => x"80",
          6835 => x"1b",
          6836 => x"db",
          6837 => x"b6",
          6838 => x"ea",
          6839 => x"98",
          6840 => x"34",
          6841 => x"51",
          6842 => x"82",
          6843 => x"83",
          6844 => x"53",
          6845 => x"d5",
          6846 => x"06",
          6847 => x"b4",
          6848 => x"84",
          6849 => x"98",
          6850 => x"85",
          6851 => x"09",
          6852 => x"38",
          6853 => x"51",
          6854 => x"82",
          6855 => x"86",
          6856 => x"f2",
          6857 => x"06",
          6858 => x"9c",
          6859 => x"d8",
          6860 => x"98",
          6861 => x"0c",
          6862 => x"51",
          6863 => x"82",
          6864 => x"8c",
          6865 => x"74",
          6866 => x"e0",
          6867 => x"53",
          6868 => x"e0",
          6869 => x"15",
          6870 => x"94",
          6871 => x"56",
          6872 => x"98",
          6873 => x"0d",
          6874 => x"0d",
          6875 => x"55",
          6876 => x"b9",
          6877 => x"53",
          6878 => x"b1",
          6879 => x"52",
          6880 => x"a9",
          6881 => x"22",
          6882 => x"57",
          6883 => x"2e",
          6884 => x"99",
          6885 => x"33",
          6886 => x"3f",
          6887 => x"08",
          6888 => x"71",
          6889 => x"74",
          6890 => x"83",
          6891 => x"78",
          6892 => x"52",
          6893 => x"98",
          6894 => x"0d",
          6895 => x"0d",
          6896 => x"33",
          6897 => x"3d",
          6898 => x"56",
          6899 => x"8b",
          6900 => x"82",
          6901 => x"24",
          6902 => x"b6",
          6903 => x"29",
          6904 => x"05",
          6905 => x"55",
          6906 => x"84",
          6907 => x"34",
          6908 => x"80",
          6909 => x"80",
          6910 => x"75",
          6911 => x"75",
          6912 => x"38",
          6913 => x"3d",
          6914 => x"05",
          6915 => x"3f",
          6916 => x"08",
          6917 => x"b6",
          6918 => x"3d",
          6919 => x"3d",
          6920 => x"84",
          6921 => x"05",
          6922 => x"89",
          6923 => x"2e",
          6924 => x"77",
          6925 => x"54",
          6926 => x"05",
          6927 => x"84",
          6928 => x"f6",
          6929 => x"b6",
          6930 => x"82",
          6931 => x"84",
          6932 => x"5c",
          6933 => x"3d",
          6934 => x"ed",
          6935 => x"b6",
          6936 => x"82",
          6937 => x"92",
          6938 => x"d7",
          6939 => x"98",
          6940 => x"73",
          6941 => x"38",
          6942 => x"9c",
          6943 => x"80",
          6944 => x"38",
          6945 => x"95",
          6946 => x"2e",
          6947 => x"aa",
          6948 => x"ea",
          6949 => x"b6",
          6950 => x"9e",
          6951 => x"05",
          6952 => x"54",
          6953 => x"38",
          6954 => x"70",
          6955 => x"54",
          6956 => x"8e",
          6957 => x"83",
          6958 => x"88",
          6959 => x"83",
          6960 => x"83",
          6961 => x"06",
          6962 => x"80",
          6963 => x"38",
          6964 => x"51",
          6965 => x"82",
          6966 => x"56",
          6967 => x"0a",
          6968 => x"05",
          6969 => x"3f",
          6970 => x"0b",
          6971 => x"80",
          6972 => x"7a",
          6973 => x"3f",
          6974 => x"9c",
          6975 => x"d1",
          6976 => x"81",
          6977 => x"34",
          6978 => x"80",
          6979 => x"b0",
          6980 => x"54",
          6981 => x"52",
          6982 => x"05",
          6983 => x"3f",
          6984 => x"08",
          6985 => x"98",
          6986 => x"38",
          6987 => x"82",
          6988 => x"b2",
          6989 => x"84",
          6990 => x"06",
          6991 => x"73",
          6992 => x"38",
          6993 => x"ad",
          6994 => x"2a",
          6995 => x"51",
          6996 => x"2e",
          6997 => x"81",
          6998 => x"80",
          6999 => x"87",
          7000 => x"39",
          7001 => x"51",
          7002 => x"82",
          7003 => x"7b",
          7004 => x"12",
          7005 => x"82",
          7006 => x"81",
          7007 => x"83",
          7008 => x"06",
          7009 => x"80",
          7010 => x"77",
          7011 => x"58",
          7012 => x"08",
          7013 => x"63",
          7014 => x"63",
          7015 => x"57",
          7016 => x"82",
          7017 => x"82",
          7018 => x"88",
          7019 => x"9c",
          7020 => x"d2",
          7021 => x"b6",
          7022 => x"b6",
          7023 => x"1b",
          7024 => x"0c",
          7025 => x"22",
          7026 => x"77",
          7027 => x"80",
          7028 => x"34",
          7029 => x"1a",
          7030 => x"94",
          7031 => x"85",
          7032 => x"06",
          7033 => x"80",
          7034 => x"38",
          7035 => x"08",
          7036 => x"84",
          7037 => x"98",
          7038 => x"0c",
          7039 => x"70",
          7040 => x"52",
          7041 => x"39",
          7042 => x"51",
          7043 => x"82",
          7044 => x"57",
          7045 => x"08",
          7046 => x"38",
          7047 => x"b6",
          7048 => x"2e",
          7049 => x"83",
          7050 => x"75",
          7051 => x"74",
          7052 => x"07",
          7053 => x"54",
          7054 => x"8a",
          7055 => x"75",
          7056 => x"73",
          7057 => x"98",
          7058 => x"a9",
          7059 => x"ff",
          7060 => x"80",
          7061 => x"76",
          7062 => x"d6",
          7063 => x"b6",
          7064 => x"38",
          7065 => x"39",
          7066 => x"82",
          7067 => x"05",
          7068 => x"84",
          7069 => x"0c",
          7070 => x"82",
          7071 => x"97",
          7072 => x"f2",
          7073 => x"63",
          7074 => x"40",
          7075 => x"7e",
          7076 => x"fc",
          7077 => x"51",
          7078 => x"82",
          7079 => x"55",
          7080 => x"08",
          7081 => x"19",
          7082 => x"80",
          7083 => x"74",
          7084 => x"39",
          7085 => x"81",
          7086 => x"56",
          7087 => x"82",
          7088 => x"39",
          7089 => x"1a",
          7090 => x"82",
          7091 => x"0b",
          7092 => x"81",
          7093 => x"39",
          7094 => x"94",
          7095 => x"55",
          7096 => x"83",
          7097 => x"7b",
          7098 => x"89",
          7099 => x"08",
          7100 => x"06",
          7101 => x"81",
          7102 => x"8a",
          7103 => x"05",
          7104 => x"06",
          7105 => x"a8",
          7106 => x"38",
          7107 => x"55",
          7108 => x"19",
          7109 => x"51",
          7110 => x"82",
          7111 => x"55",
          7112 => x"ff",
          7113 => x"ff",
          7114 => x"38",
          7115 => x"0c",
          7116 => x"52",
          7117 => x"cb",
          7118 => x"98",
          7119 => x"ff",
          7120 => x"b6",
          7121 => x"7c",
          7122 => x"57",
          7123 => x"80",
          7124 => x"1a",
          7125 => x"22",
          7126 => x"75",
          7127 => x"38",
          7128 => x"58",
          7129 => x"53",
          7130 => x"1b",
          7131 => x"88",
          7132 => x"98",
          7133 => x"38",
          7134 => x"33",
          7135 => x"80",
          7136 => x"b0",
          7137 => x"31",
          7138 => x"27",
          7139 => x"80",
          7140 => x"52",
          7141 => x"77",
          7142 => x"7d",
          7143 => x"e0",
          7144 => x"2b",
          7145 => x"76",
          7146 => x"94",
          7147 => x"ff",
          7148 => x"71",
          7149 => x"7b",
          7150 => x"38",
          7151 => x"19",
          7152 => x"51",
          7153 => x"82",
          7154 => x"fe",
          7155 => x"53",
          7156 => x"83",
          7157 => x"b4",
          7158 => x"51",
          7159 => x"7b",
          7160 => x"08",
          7161 => x"76",
          7162 => x"08",
          7163 => x"0c",
          7164 => x"f3",
          7165 => x"75",
          7166 => x"0c",
          7167 => x"04",
          7168 => x"60",
          7169 => x"40",
          7170 => x"80",
          7171 => x"3d",
          7172 => x"77",
          7173 => x"3f",
          7174 => x"08",
          7175 => x"98",
          7176 => x"91",
          7177 => x"74",
          7178 => x"38",
          7179 => x"b8",
          7180 => x"33",
          7181 => x"70",
          7182 => x"56",
          7183 => x"74",
          7184 => x"a4",
          7185 => x"82",
          7186 => x"34",
          7187 => x"98",
          7188 => x"91",
          7189 => x"56",
          7190 => x"94",
          7191 => x"11",
          7192 => x"76",
          7193 => x"75",
          7194 => x"80",
          7195 => x"38",
          7196 => x"70",
          7197 => x"56",
          7198 => x"fd",
          7199 => x"11",
          7200 => x"77",
          7201 => x"5c",
          7202 => x"38",
          7203 => x"88",
          7204 => x"74",
          7205 => x"52",
          7206 => x"18",
          7207 => x"51",
          7208 => x"82",
          7209 => x"55",
          7210 => x"08",
          7211 => x"ab",
          7212 => x"2e",
          7213 => x"74",
          7214 => x"95",
          7215 => x"19",
          7216 => x"08",
          7217 => x"88",
          7218 => x"55",
          7219 => x"9c",
          7220 => x"09",
          7221 => x"38",
          7222 => x"c1",
          7223 => x"98",
          7224 => x"38",
          7225 => x"52",
          7226 => x"97",
          7227 => x"98",
          7228 => x"fe",
          7229 => x"b6",
          7230 => x"7c",
          7231 => x"57",
          7232 => x"80",
          7233 => x"1b",
          7234 => x"22",
          7235 => x"75",
          7236 => x"38",
          7237 => x"59",
          7238 => x"53",
          7239 => x"1a",
          7240 => x"be",
          7241 => x"98",
          7242 => x"38",
          7243 => x"08",
          7244 => x"56",
          7245 => x"9b",
          7246 => x"53",
          7247 => x"77",
          7248 => x"7d",
          7249 => x"16",
          7250 => x"3f",
          7251 => x"0b",
          7252 => x"78",
          7253 => x"80",
          7254 => x"18",
          7255 => x"08",
          7256 => x"7e",
          7257 => x"3f",
          7258 => x"08",
          7259 => x"7e",
          7260 => x"0c",
          7261 => x"19",
          7262 => x"08",
          7263 => x"84",
          7264 => x"57",
          7265 => x"27",
          7266 => x"56",
          7267 => x"52",
          7268 => x"f9",
          7269 => x"98",
          7270 => x"38",
          7271 => x"52",
          7272 => x"83",
          7273 => x"b4",
          7274 => x"d4",
          7275 => x"81",
          7276 => x"34",
          7277 => x"7e",
          7278 => x"0c",
          7279 => x"1a",
          7280 => x"94",
          7281 => x"1b",
          7282 => x"5e",
          7283 => x"27",
          7284 => x"55",
          7285 => x"0c",
          7286 => x"90",
          7287 => x"c0",
          7288 => x"90",
          7289 => x"56",
          7290 => x"98",
          7291 => x"0d",
          7292 => x"0d",
          7293 => x"fc",
          7294 => x"52",
          7295 => x"3f",
          7296 => x"08",
          7297 => x"98",
          7298 => x"38",
          7299 => x"70",
          7300 => x"81",
          7301 => x"55",
          7302 => x"80",
          7303 => x"16",
          7304 => x"51",
          7305 => x"82",
          7306 => x"57",
          7307 => x"08",
          7308 => x"a4",
          7309 => x"11",
          7310 => x"55",
          7311 => x"16",
          7312 => x"08",
          7313 => x"75",
          7314 => x"e8",
          7315 => x"08",
          7316 => x"51",
          7317 => x"82",
          7318 => x"52",
          7319 => x"c9",
          7320 => x"52",
          7321 => x"c9",
          7322 => x"54",
          7323 => x"15",
          7324 => x"cc",
          7325 => x"b6",
          7326 => x"17",
          7327 => x"06",
          7328 => x"90",
          7329 => x"82",
          7330 => x"8a",
          7331 => x"fc",
          7332 => x"70",
          7333 => x"d9",
          7334 => x"98",
          7335 => x"b6",
          7336 => x"38",
          7337 => x"05",
          7338 => x"f1",
          7339 => x"b6",
          7340 => x"82",
          7341 => x"87",
          7342 => x"98",
          7343 => x"72",
          7344 => x"0c",
          7345 => x"04",
          7346 => x"84",
          7347 => x"e4",
          7348 => x"80",
          7349 => x"98",
          7350 => x"38",
          7351 => x"08",
          7352 => x"34",
          7353 => x"82",
          7354 => x"83",
          7355 => x"ef",
          7356 => x"53",
          7357 => x"05",
          7358 => x"51",
          7359 => x"82",
          7360 => x"55",
          7361 => x"08",
          7362 => x"76",
          7363 => x"93",
          7364 => x"51",
          7365 => x"82",
          7366 => x"55",
          7367 => x"08",
          7368 => x"80",
          7369 => x"70",
          7370 => x"56",
          7371 => x"89",
          7372 => x"94",
          7373 => x"b2",
          7374 => x"05",
          7375 => x"2a",
          7376 => x"51",
          7377 => x"80",
          7378 => x"76",
          7379 => x"52",
          7380 => x"3f",
          7381 => x"08",
          7382 => x"8e",
          7383 => x"98",
          7384 => x"09",
          7385 => x"38",
          7386 => x"82",
          7387 => x"93",
          7388 => x"e4",
          7389 => x"6f",
          7390 => x"7a",
          7391 => x"9e",
          7392 => x"05",
          7393 => x"51",
          7394 => x"82",
          7395 => x"57",
          7396 => x"08",
          7397 => x"7b",
          7398 => x"94",
          7399 => x"55",
          7400 => x"73",
          7401 => x"ed",
          7402 => x"93",
          7403 => x"55",
          7404 => x"82",
          7405 => x"57",
          7406 => x"08",
          7407 => x"68",
          7408 => x"c9",
          7409 => x"b6",
          7410 => x"82",
          7411 => x"82",
          7412 => x"52",
          7413 => x"a3",
          7414 => x"98",
          7415 => x"52",
          7416 => x"b8",
          7417 => x"98",
          7418 => x"b6",
          7419 => x"a2",
          7420 => x"74",
          7421 => x"3f",
          7422 => x"08",
          7423 => x"98",
          7424 => x"69",
          7425 => x"d9",
          7426 => x"82",
          7427 => x"2e",
          7428 => x"52",
          7429 => x"cf",
          7430 => x"98",
          7431 => x"b6",
          7432 => x"2e",
          7433 => x"84",
          7434 => x"06",
          7435 => x"57",
          7436 => x"76",
          7437 => x"9e",
          7438 => x"05",
          7439 => x"dc",
          7440 => x"90",
          7441 => x"81",
          7442 => x"56",
          7443 => x"80",
          7444 => x"02",
          7445 => x"81",
          7446 => x"70",
          7447 => x"56",
          7448 => x"81",
          7449 => x"78",
          7450 => x"38",
          7451 => x"99",
          7452 => x"81",
          7453 => x"18",
          7454 => x"18",
          7455 => x"58",
          7456 => x"33",
          7457 => x"ee",
          7458 => x"6f",
          7459 => x"af",
          7460 => x"8d",
          7461 => x"2e",
          7462 => x"8a",
          7463 => x"6f",
          7464 => x"af",
          7465 => x"0b",
          7466 => x"33",
          7467 => x"82",
          7468 => x"70",
          7469 => x"52",
          7470 => x"56",
          7471 => x"8d",
          7472 => x"70",
          7473 => x"51",
          7474 => x"f5",
          7475 => x"54",
          7476 => x"a7",
          7477 => x"74",
          7478 => x"38",
          7479 => x"73",
          7480 => x"81",
          7481 => x"81",
          7482 => x"39",
          7483 => x"81",
          7484 => x"74",
          7485 => x"81",
          7486 => x"91",
          7487 => x"6e",
          7488 => x"59",
          7489 => x"7a",
          7490 => x"5c",
          7491 => x"26",
          7492 => x"7a",
          7493 => x"b6",
          7494 => x"3d",
          7495 => x"3d",
          7496 => x"8d",
          7497 => x"54",
          7498 => x"55",
          7499 => x"82",
          7500 => x"53",
          7501 => x"08",
          7502 => x"91",
          7503 => x"72",
          7504 => x"8c",
          7505 => x"73",
          7506 => x"38",
          7507 => x"70",
          7508 => x"81",
          7509 => x"57",
          7510 => x"73",
          7511 => x"08",
          7512 => x"94",
          7513 => x"75",
          7514 => x"97",
          7515 => x"11",
          7516 => x"2b",
          7517 => x"73",
          7518 => x"38",
          7519 => x"16",
          7520 => x"ff",
          7521 => x"98",
          7522 => x"78",
          7523 => x"55",
          7524 => x"ef",
          7525 => x"98",
          7526 => x"96",
          7527 => x"70",
          7528 => x"94",
          7529 => x"71",
          7530 => x"08",
          7531 => x"53",
          7532 => x"15",
          7533 => x"a6",
          7534 => x"74",
          7535 => x"3f",
          7536 => x"08",
          7537 => x"98",
          7538 => x"81",
          7539 => x"b6",
          7540 => x"2e",
          7541 => x"82",
          7542 => x"88",
          7543 => x"98",
          7544 => x"80",
          7545 => x"38",
          7546 => x"80",
          7547 => x"77",
          7548 => x"08",
          7549 => x"0c",
          7550 => x"70",
          7551 => x"81",
          7552 => x"5a",
          7553 => x"2e",
          7554 => x"52",
          7555 => x"f9",
          7556 => x"98",
          7557 => x"b6",
          7558 => x"38",
          7559 => x"08",
          7560 => x"73",
          7561 => x"c7",
          7562 => x"b6",
          7563 => x"73",
          7564 => x"38",
          7565 => x"af",
          7566 => x"73",
          7567 => x"27",
          7568 => x"98",
          7569 => x"a0",
          7570 => x"08",
          7571 => x"0c",
          7572 => x"06",
          7573 => x"2e",
          7574 => x"52",
          7575 => x"a3",
          7576 => x"98",
          7577 => x"82",
          7578 => x"34",
          7579 => x"c4",
          7580 => x"91",
          7581 => x"53",
          7582 => x"89",
          7583 => x"98",
          7584 => x"94",
          7585 => x"8c",
          7586 => x"27",
          7587 => x"8c",
          7588 => x"15",
          7589 => x"07",
          7590 => x"16",
          7591 => x"ff",
          7592 => x"80",
          7593 => x"77",
          7594 => x"2e",
          7595 => x"9c",
          7596 => x"53",
          7597 => x"98",
          7598 => x"0d",
          7599 => x"0d",
          7600 => x"54",
          7601 => x"81",
          7602 => x"53",
          7603 => x"05",
          7604 => x"84",
          7605 => x"e7",
          7606 => x"98",
          7607 => x"b6",
          7608 => x"ea",
          7609 => x"0c",
          7610 => x"51",
          7611 => x"82",
          7612 => x"55",
          7613 => x"08",
          7614 => x"ab",
          7615 => x"98",
          7616 => x"80",
          7617 => x"38",
          7618 => x"70",
          7619 => x"81",
          7620 => x"57",
          7621 => x"ad",
          7622 => x"08",
          7623 => x"d3",
          7624 => x"b6",
          7625 => x"17",
          7626 => x"86",
          7627 => x"17",
          7628 => x"75",
          7629 => x"3f",
          7630 => x"08",
          7631 => x"2e",
          7632 => x"85",
          7633 => x"86",
          7634 => x"2e",
          7635 => x"76",
          7636 => x"73",
          7637 => x"0c",
          7638 => x"04",
          7639 => x"76",
          7640 => x"05",
          7641 => x"53",
          7642 => x"82",
          7643 => x"87",
          7644 => x"98",
          7645 => x"86",
          7646 => x"fb",
          7647 => x"79",
          7648 => x"05",
          7649 => x"56",
          7650 => x"3f",
          7651 => x"08",
          7652 => x"98",
          7653 => x"38",
          7654 => x"82",
          7655 => x"52",
          7656 => x"f8",
          7657 => x"98",
          7658 => x"ca",
          7659 => x"98",
          7660 => x"51",
          7661 => x"82",
          7662 => x"53",
          7663 => x"08",
          7664 => x"81",
          7665 => x"80",
          7666 => x"82",
          7667 => x"a6",
          7668 => x"73",
          7669 => x"3f",
          7670 => x"51",
          7671 => x"82",
          7672 => x"84",
          7673 => x"70",
          7674 => x"2c",
          7675 => x"98",
          7676 => x"51",
          7677 => x"82",
          7678 => x"87",
          7679 => x"ee",
          7680 => x"57",
          7681 => x"3d",
          7682 => x"3d",
          7683 => x"af",
          7684 => x"98",
          7685 => x"b6",
          7686 => x"38",
          7687 => x"51",
          7688 => x"82",
          7689 => x"55",
          7690 => x"08",
          7691 => x"80",
          7692 => x"70",
          7693 => x"58",
          7694 => x"85",
          7695 => x"8d",
          7696 => x"2e",
          7697 => x"52",
          7698 => x"be",
          7699 => x"b6",
          7700 => x"3d",
          7701 => x"3d",
          7702 => x"55",
          7703 => x"92",
          7704 => x"52",
          7705 => x"de",
          7706 => x"b6",
          7707 => x"82",
          7708 => x"82",
          7709 => x"74",
          7710 => x"98",
          7711 => x"11",
          7712 => x"59",
          7713 => x"75",
          7714 => x"38",
          7715 => x"81",
          7716 => x"5b",
          7717 => x"82",
          7718 => x"39",
          7719 => x"08",
          7720 => x"59",
          7721 => x"09",
          7722 => x"38",
          7723 => x"57",
          7724 => x"3d",
          7725 => x"c1",
          7726 => x"b6",
          7727 => x"2e",
          7728 => x"b6",
          7729 => x"2e",
          7730 => x"b6",
          7731 => x"70",
          7732 => x"08",
          7733 => x"7a",
          7734 => x"7f",
          7735 => x"54",
          7736 => x"77",
          7737 => x"80",
          7738 => x"15",
          7739 => x"98",
          7740 => x"75",
          7741 => x"52",
          7742 => x"52",
          7743 => x"8d",
          7744 => x"98",
          7745 => x"b6",
          7746 => x"d6",
          7747 => x"33",
          7748 => x"1a",
          7749 => x"54",
          7750 => x"09",
          7751 => x"38",
          7752 => x"ff",
          7753 => x"82",
          7754 => x"83",
          7755 => x"70",
          7756 => x"25",
          7757 => x"59",
          7758 => x"9b",
          7759 => x"51",
          7760 => x"3f",
          7761 => x"08",
          7762 => x"70",
          7763 => x"25",
          7764 => x"59",
          7765 => x"75",
          7766 => x"7a",
          7767 => x"ff",
          7768 => x"7c",
          7769 => x"90",
          7770 => x"11",
          7771 => x"56",
          7772 => x"15",
          7773 => x"b6",
          7774 => x"3d",
          7775 => x"3d",
          7776 => x"3d",
          7777 => x"70",
          7778 => x"dd",
          7779 => x"98",
          7780 => x"b6",
          7781 => x"a8",
          7782 => x"33",
          7783 => x"a0",
          7784 => x"33",
          7785 => x"70",
          7786 => x"55",
          7787 => x"73",
          7788 => x"8e",
          7789 => x"08",
          7790 => x"18",
          7791 => x"80",
          7792 => x"38",
          7793 => x"08",
          7794 => x"08",
          7795 => x"c4",
          7796 => x"b6",
          7797 => x"88",
          7798 => x"80",
          7799 => x"17",
          7800 => x"51",
          7801 => x"3f",
          7802 => x"08",
          7803 => x"81",
          7804 => x"81",
          7805 => x"98",
          7806 => x"09",
          7807 => x"38",
          7808 => x"39",
          7809 => x"77",
          7810 => x"98",
          7811 => x"08",
          7812 => x"98",
          7813 => x"82",
          7814 => x"52",
          7815 => x"bd",
          7816 => x"98",
          7817 => x"17",
          7818 => x"0c",
          7819 => x"80",
          7820 => x"73",
          7821 => x"75",
          7822 => x"38",
          7823 => x"34",
          7824 => x"82",
          7825 => x"89",
          7826 => x"e2",
          7827 => x"53",
          7828 => x"a4",
          7829 => x"3d",
          7830 => x"3f",
          7831 => x"08",
          7832 => x"98",
          7833 => x"38",
          7834 => x"3d",
          7835 => x"3d",
          7836 => x"d1",
          7837 => x"b6",
          7838 => x"82",
          7839 => x"81",
          7840 => x"80",
          7841 => x"70",
          7842 => x"81",
          7843 => x"56",
          7844 => x"81",
          7845 => x"98",
          7846 => x"74",
          7847 => x"38",
          7848 => x"05",
          7849 => x"06",
          7850 => x"55",
          7851 => x"38",
          7852 => x"51",
          7853 => x"82",
          7854 => x"74",
          7855 => x"81",
          7856 => x"56",
          7857 => x"80",
          7858 => x"54",
          7859 => x"08",
          7860 => x"2e",
          7861 => x"73",
          7862 => x"98",
          7863 => x"52",
          7864 => x"52",
          7865 => x"3f",
          7866 => x"08",
          7867 => x"98",
          7868 => x"38",
          7869 => x"08",
          7870 => x"cc",
          7871 => x"b6",
          7872 => x"82",
          7873 => x"86",
          7874 => x"80",
          7875 => x"b6",
          7876 => x"2e",
          7877 => x"b6",
          7878 => x"c0",
          7879 => x"ce",
          7880 => x"b6",
          7881 => x"b6",
          7882 => x"70",
          7883 => x"08",
          7884 => x"51",
          7885 => x"80",
          7886 => x"73",
          7887 => x"38",
          7888 => x"52",
          7889 => x"95",
          7890 => x"98",
          7891 => x"8c",
          7892 => x"ff",
          7893 => x"82",
          7894 => x"55",
          7895 => x"98",
          7896 => x"0d",
          7897 => x"0d",
          7898 => x"3d",
          7899 => x"9a",
          7900 => x"cb",
          7901 => x"98",
          7902 => x"b6",
          7903 => x"b0",
          7904 => x"69",
          7905 => x"70",
          7906 => x"97",
          7907 => x"98",
          7908 => x"b6",
          7909 => x"38",
          7910 => x"94",
          7911 => x"98",
          7912 => x"09",
          7913 => x"88",
          7914 => x"df",
          7915 => x"85",
          7916 => x"51",
          7917 => x"74",
          7918 => x"78",
          7919 => x"8a",
          7920 => x"57",
          7921 => x"82",
          7922 => x"75",
          7923 => x"b6",
          7924 => x"38",
          7925 => x"b6",
          7926 => x"2e",
          7927 => x"83",
          7928 => x"82",
          7929 => x"ff",
          7930 => x"06",
          7931 => x"54",
          7932 => x"73",
          7933 => x"82",
          7934 => x"52",
          7935 => x"a4",
          7936 => x"98",
          7937 => x"b6",
          7938 => x"9a",
          7939 => x"a0",
          7940 => x"51",
          7941 => x"3f",
          7942 => x"0b",
          7943 => x"78",
          7944 => x"bf",
          7945 => x"88",
          7946 => x"80",
          7947 => x"ff",
          7948 => x"75",
          7949 => x"11",
          7950 => x"f8",
          7951 => x"78",
          7952 => x"80",
          7953 => x"ff",
          7954 => x"78",
          7955 => x"80",
          7956 => x"7f",
          7957 => x"d4",
          7958 => x"c9",
          7959 => x"54",
          7960 => x"15",
          7961 => x"cb",
          7962 => x"b6",
          7963 => x"82",
          7964 => x"b2",
          7965 => x"b2",
          7966 => x"96",
          7967 => x"b5",
          7968 => x"53",
          7969 => x"51",
          7970 => x"64",
          7971 => x"8b",
          7972 => x"54",
          7973 => x"15",
          7974 => x"ff",
          7975 => x"82",
          7976 => x"54",
          7977 => x"53",
          7978 => x"51",
          7979 => x"3f",
          7980 => x"98",
          7981 => x"0d",
          7982 => x"0d",
          7983 => x"05",
          7984 => x"3f",
          7985 => x"3d",
          7986 => x"52",
          7987 => x"d5",
          7988 => x"b6",
          7989 => x"82",
          7990 => x"82",
          7991 => x"4d",
          7992 => x"52",
          7993 => x"52",
          7994 => x"3f",
          7995 => x"08",
          7996 => x"98",
          7997 => x"38",
          7998 => x"05",
          7999 => x"06",
          8000 => x"73",
          8001 => x"a0",
          8002 => x"08",
          8003 => x"ff",
          8004 => x"ff",
          8005 => x"ac",
          8006 => x"92",
          8007 => x"54",
          8008 => x"3f",
          8009 => x"52",
          8010 => x"f7",
          8011 => x"98",
          8012 => x"b6",
          8013 => x"38",
          8014 => x"09",
          8015 => x"38",
          8016 => x"08",
          8017 => x"88",
          8018 => x"39",
          8019 => x"08",
          8020 => x"81",
          8021 => x"38",
          8022 => x"b1",
          8023 => x"98",
          8024 => x"b6",
          8025 => x"c8",
          8026 => x"93",
          8027 => x"ff",
          8028 => x"8d",
          8029 => x"b4",
          8030 => x"af",
          8031 => x"17",
          8032 => x"33",
          8033 => x"70",
          8034 => x"55",
          8035 => x"38",
          8036 => x"54",
          8037 => x"34",
          8038 => x"0b",
          8039 => x"8b",
          8040 => x"84",
          8041 => x"06",
          8042 => x"73",
          8043 => x"e5",
          8044 => x"2e",
          8045 => x"75",
          8046 => x"c6",
          8047 => x"b6",
          8048 => x"78",
          8049 => x"bb",
          8050 => x"82",
          8051 => x"80",
          8052 => x"38",
          8053 => x"08",
          8054 => x"ff",
          8055 => x"82",
          8056 => x"79",
          8057 => x"58",
          8058 => x"b6",
          8059 => x"c0",
          8060 => x"33",
          8061 => x"2e",
          8062 => x"99",
          8063 => x"75",
          8064 => x"c6",
          8065 => x"54",
          8066 => x"15",
          8067 => x"82",
          8068 => x"9c",
          8069 => x"c8",
          8070 => x"b6",
          8071 => x"82",
          8072 => x"8c",
          8073 => x"ff",
          8074 => x"82",
          8075 => x"55",
          8076 => x"98",
          8077 => x"0d",
          8078 => x"0d",
          8079 => x"05",
          8080 => x"05",
          8081 => x"33",
          8082 => x"53",
          8083 => x"05",
          8084 => x"51",
          8085 => x"82",
          8086 => x"55",
          8087 => x"08",
          8088 => x"78",
          8089 => x"95",
          8090 => x"51",
          8091 => x"82",
          8092 => x"55",
          8093 => x"08",
          8094 => x"80",
          8095 => x"81",
          8096 => x"86",
          8097 => x"38",
          8098 => x"61",
          8099 => x"12",
          8100 => x"7a",
          8101 => x"51",
          8102 => x"74",
          8103 => x"78",
          8104 => x"83",
          8105 => x"51",
          8106 => x"3f",
          8107 => x"08",
          8108 => x"b6",
          8109 => x"3d",
          8110 => x"3d",
          8111 => x"82",
          8112 => x"d0",
          8113 => x"3d",
          8114 => x"3f",
          8115 => x"08",
          8116 => x"98",
          8117 => x"38",
          8118 => x"52",
          8119 => x"05",
          8120 => x"3f",
          8121 => x"08",
          8122 => x"98",
          8123 => x"02",
          8124 => x"33",
          8125 => x"54",
          8126 => x"a6",
          8127 => x"22",
          8128 => x"71",
          8129 => x"53",
          8130 => x"51",
          8131 => x"3f",
          8132 => x"0b",
          8133 => x"76",
          8134 => x"b8",
          8135 => x"98",
          8136 => x"82",
          8137 => x"93",
          8138 => x"ea",
          8139 => x"6b",
          8140 => x"53",
          8141 => x"05",
          8142 => x"51",
          8143 => x"82",
          8144 => x"82",
          8145 => x"30",
          8146 => x"98",
          8147 => x"25",
          8148 => x"79",
          8149 => x"85",
          8150 => x"75",
          8151 => x"73",
          8152 => x"f9",
          8153 => x"80",
          8154 => x"8d",
          8155 => x"54",
          8156 => x"3f",
          8157 => x"08",
          8158 => x"98",
          8159 => x"38",
          8160 => x"51",
          8161 => x"82",
          8162 => x"57",
          8163 => x"08",
          8164 => x"b6",
          8165 => x"b6",
          8166 => x"5b",
          8167 => x"18",
          8168 => x"18",
          8169 => x"74",
          8170 => x"81",
          8171 => x"78",
          8172 => x"8b",
          8173 => x"54",
          8174 => x"75",
          8175 => x"38",
          8176 => x"1b",
          8177 => x"55",
          8178 => x"2e",
          8179 => x"39",
          8180 => x"09",
          8181 => x"38",
          8182 => x"80",
          8183 => x"70",
          8184 => x"25",
          8185 => x"80",
          8186 => x"38",
          8187 => x"bc",
          8188 => x"11",
          8189 => x"ff",
          8190 => x"82",
          8191 => x"57",
          8192 => x"08",
          8193 => x"70",
          8194 => x"80",
          8195 => x"83",
          8196 => x"80",
          8197 => x"84",
          8198 => x"a7",
          8199 => x"b4",
          8200 => x"ad",
          8201 => x"b6",
          8202 => x"0c",
          8203 => x"98",
          8204 => x"0d",
          8205 => x"0d",
          8206 => x"3d",
          8207 => x"52",
          8208 => x"ce",
          8209 => x"b6",
          8210 => x"b6",
          8211 => x"54",
          8212 => x"08",
          8213 => x"8b",
          8214 => x"8b",
          8215 => x"59",
          8216 => x"3f",
          8217 => x"33",
          8218 => x"06",
          8219 => x"57",
          8220 => x"81",
          8221 => x"58",
          8222 => x"06",
          8223 => x"4e",
          8224 => x"ff",
          8225 => x"82",
          8226 => x"80",
          8227 => x"6c",
          8228 => x"53",
          8229 => x"ae",
          8230 => x"b6",
          8231 => x"2e",
          8232 => x"88",
          8233 => x"6d",
          8234 => x"55",
          8235 => x"b6",
          8236 => x"ff",
          8237 => x"83",
          8238 => x"51",
          8239 => x"26",
          8240 => x"15",
          8241 => x"ff",
          8242 => x"80",
          8243 => x"87",
          8244 => x"e0",
          8245 => x"74",
          8246 => x"38",
          8247 => x"b0",
          8248 => x"ae",
          8249 => x"b6",
          8250 => x"38",
          8251 => x"27",
          8252 => x"89",
          8253 => x"8b",
          8254 => x"27",
          8255 => x"55",
          8256 => x"81",
          8257 => x"8f",
          8258 => x"2a",
          8259 => x"70",
          8260 => x"34",
          8261 => x"74",
          8262 => x"05",
          8263 => x"17",
          8264 => x"70",
          8265 => x"52",
          8266 => x"73",
          8267 => x"c8",
          8268 => x"33",
          8269 => x"73",
          8270 => x"81",
          8271 => x"80",
          8272 => x"02",
          8273 => x"76",
          8274 => x"51",
          8275 => x"2e",
          8276 => x"87",
          8277 => x"57",
          8278 => x"79",
          8279 => x"80",
          8280 => x"70",
          8281 => x"ba",
          8282 => x"b6",
          8283 => x"82",
          8284 => x"80",
          8285 => x"52",
          8286 => x"bf",
          8287 => x"b6",
          8288 => x"82",
          8289 => x"8d",
          8290 => x"c4",
          8291 => x"e5",
          8292 => x"c6",
          8293 => x"98",
          8294 => x"09",
          8295 => x"cc",
          8296 => x"76",
          8297 => x"c4",
          8298 => x"74",
          8299 => x"b0",
          8300 => x"98",
          8301 => x"b6",
          8302 => x"38",
          8303 => x"b6",
          8304 => x"67",
          8305 => x"db",
          8306 => x"88",
          8307 => x"34",
          8308 => x"52",
          8309 => x"ab",
          8310 => x"54",
          8311 => x"15",
          8312 => x"ff",
          8313 => x"82",
          8314 => x"54",
          8315 => x"82",
          8316 => x"9c",
          8317 => x"f2",
          8318 => x"62",
          8319 => x"80",
          8320 => x"93",
          8321 => x"55",
          8322 => x"5e",
          8323 => x"3f",
          8324 => x"08",
          8325 => x"98",
          8326 => x"38",
          8327 => x"58",
          8328 => x"38",
          8329 => x"97",
          8330 => x"08",
          8331 => x"38",
          8332 => x"70",
          8333 => x"81",
          8334 => x"55",
          8335 => x"87",
          8336 => x"39",
          8337 => x"90",
          8338 => x"82",
          8339 => x"8a",
          8340 => x"89",
          8341 => x"7f",
          8342 => x"56",
          8343 => x"3f",
          8344 => x"06",
          8345 => x"72",
          8346 => x"82",
          8347 => x"05",
          8348 => x"7c",
          8349 => x"55",
          8350 => x"27",
          8351 => x"16",
          8352 => x"83",
          8353 => x"76",
          8354 => x"80",
          8355 => x"79",
          8356 => x"99",
          8357 => x"7f",
          8358 => x"14",
          8359 => x"83",
          8360 => x"82",
          8361 => x"81",
          8362 => x"38",
          8363 => x"08",
          8364 => x"95",
          8365 => x"98",
          8366 => x"81",
          8367 => x"7b",
          8368 => x"06",
          8369 => x"39",
          8370 => x"56",
          8371 => x"09",
          8372 => x"b9",
          8373 => x"80",
          8374 => x"80",
          8375 => x"78",
          8376 => x"7a",
          8377 => x"38",
          8378 => x"73",
          8379 => x"81",
          8380 => x"ff",
          8381 => x"74",
          8382 => x"ff",
          8383 => x"82",
          8384 => x"58",
          8385 => x"08",
          8386 => x"74",
          8387 => x"16",
          8388 => x"73",
          8389 => x"39",
          8390 => x"7e",
          8391 => x"0c",
          8392 => x"2e",
          8393 => x"88",
          8394 => x"8c",
          8395 => x"1a",
          8396 => x"07",
          8397 => x"1b",
          8398 => x"08",
          8399 => x"16",
          8400 => x"75",
          8401 => x"38",
          8402 => x"90",
          8403 => x"15",
          8404 => x"54",
          8405 => x"34",
          8406 => x"82",
          8407 => x"90",
          8408 => x"e9",
          8409 => x"6d",
          8410 => x"80",
          8411 => x"9d",
          8412 => x"5c",
          8413 => x"3f",
          8414 => x"0b",
          8415 => x"08",
          8416 => x"38",
          8417 => x"08",
          8418 => x"cd",
          8419 => x"08",
          8420 => x"80",
          8421 => x"80",
          8422 => x"b6",
          8423 => x"ff",
          8424 => x"52",
          8425 => x"a0",
          8426 => x"b6",
          8427 => x"ff",
          8428 => x"06",
          8429 => x"56",
          8430 => x"38",
          8431 => x"70",
          8432 => x"55",
          8433 => x"8b",
          8434 => x"3d",
          8435 => x"83",
          8436 => x"ff",
          8437 => x"82",
          8438 => x"99",
          8439 => x"74",
          8440 => x"38",
          8441 => x"80",
          8442 => x"ff",
          8443 => x"55",
          8444 => x"83",
          8445 => x"78",
          8446 => x"38",
          8447 => x"26",
          8448 => x"81",
          8449 => x"8b",
          8450 => x"79",
          8451 => x"80",
          8452 => x"93",
          8453 => x"39",
          8454 => x"6e",
          8455 => x"89",
          8456 => x"48",
          8457 => x"83",
          8458 => x"61",
          8459 => x"25",
          8460 => x"55",
          8461 => x"8a",
          8462 => x"3d",
          8463 => x"81",
          8464 => x"ff",
          8465 => x"81",
          8466 => x"98",
          8467 => x"38",
          8468 => x"70",
          8469 => x"b6",
          8470 => x"56",
          8471 => x"38",
          8472 => x"55",
          8473 => x"75",
          8474 => x"38",
          8475 => x"70",
          8476 => x"ff",
          8477 => x"83",
          8478 => x"78",
          8479 => x"89",
          8480 => x"81",
          8481 => x"06",
          8482 => x"80",
          8483 => x"77",
          8484 => x"74",
          8485 => x"8d",
          8486 => x"06",
          8487 => x"2e",
          8488 => x"77",
          8489 => x"93",
          8490 => x"74",
          8491 => x"cb",
          8492 => x"7d",
          8493 => x"81",
          8494 => x"38",
          8495 => x"66",
          8496 => x"81",
          8497 => x"84",
          8498 => x"74",
          8499 => x"38",
          8500 => x"98",
          8501 => x"84",
          8502 => x"82",
          8503 => x"57",
          8504 => x"80",
          8505 => x"76",
          8506 => x"38",
          8507 => x"51",
          8508 => x"3f",
          8509 => x"08",
          8510 => x"87",
          8511 => x"2a",
          8512 => x"5c",
          8513 => x"b6",
          8514 => x"80",
          8515 => x"44",
          8516 => x"0a",
          8517 => x"ec",
          8518 => x"39",
          8519 => x"66",
          8520 => x"81",
          8521 => x"f4",
          8522 => x"74",
          8523 => x"38",
          8524 => x"98",
          8525 => x"f4",
          8526 => x"82",
          8527 => x"57",
          8528 => x"80",
          8529 => x"76",
          8530 => x"38",
          8531 => x"51",
          8532 => x"3f",
          8533 => x"08",
          8534 => x"57",
          8535 => x"08",
          8536 => x"96",
          8537 => x"82",
          8538 => x"10",
          8539 => x"08",
          8540 => x"72",
          8541 => x"59",
          8542 => x"ff",
          8543 => x"5d",
          8544 => x"44",
          8545 => x"11",
          8546 => x"70",
          8547 => x"71",
          8548 => x"06",
          8549 => x"52",
          8550 => x"40",
          8551 => x"09",
          8552 => x"38",
          8553 => x"18",
          8554 => x"39",
          8555 => x"79",
          8556 => x"70",
          8557 => x"58",
          8558 => x"76",
          8559 => x"38",
          8560 => x"7d",
          8561 => x"70",
          8562 => x"55",
          8563 => x"3f",
          8564 => x"08",
          8565 => x"2e",
          8566 => x"9b",
          8567 => x"98",
          8568 => x"f5",
          8569 => x"38",
          8570 => x"38",
          8571 => x"59",
          8572 => x"38",
          8573 => x"7d",
          8574 => x"81",
          8575 => x"38",
          8576 => x"0b",
          8577 => x"08",
          8578 => x"78",
          8579 => x"1a",
          8580 => x"c0",
          8581 => x"74",
          8582 => x"39",
          8583 => x"55",
          8584 => x"8f",
          8585 => x"fd",
          8586 => x"b6",
          8587 => x"f5",
          8588 => x"78",
          8589 => x"79",
          8590 => x"80",
          8591 => x"f1",
          8592 => x"39",
          8593 => x"81",
          8594 => x"06",
          8595 => x"55",
          8596 => x"27",
          8597 => x"81",
          8598 => x"56",
          8599 => x"38",
          8600 => x"80",
          8601 => x"ff",
          8602 => x"8b",
          8603 => x"9c",
          8604 => x"ff",
          8605 => x"84",
          8606 => x"1b",
          8607 => x"b3",
          8608 => x"1c",
          8609 => x"ff",
          8610 => x"8e",
          8611 => x"a1",
          8612 => x"0b",
          8613 => x"7d",
          8614 => x"30",
          8615 => x"84",
          8616 => x"51",
          8617 => x"51",
          8618 => x"3f",
          8619 => x"83",
          8620 => x"90",
          8621 => x"ff",
          8622 => x"93",
          8623 => x"a0",
          8624 => x"39",
          8625 => x"1b",
          8626 => x"85",
          8627 => x"95",
          8628 => x"52",
          8629 => x"ff",
          8630 => x"81",
          8631 => x"1b",
          8632 => x"cf",
          8633 => x"9c",
          8634 => x"a0",
          8635 => x"83",
          8636 => x"06",
          8637 => x"82",
          8638 => x"52",
          8639 => x"51",
          8640 => x"3f",
          8641 => x"1b",
          8642 => x"c5",
          8643 => x"ac",
          8644 => x"a0",
          8645 => x"52",
          8646 => x"ff",
          8647 => x"86",
          8648 => x"51",
          8649 => x"3f",
          8650 => x"80",
          8651 => x"a9",
          8652 => x"1c",
          8653 => x"82",
          8654 => x"80",
          8655 => x"ae",
          8656 => x"b2",
          8657 => x"1b",
          8658 => x"85",
          8659 => x"ff",
          8660 => x"96",
          8661 => x"9f",
          8662 => x"80",
          8663 => x"34",
          8664 => x"1c",
          8665 => x"82",
          8666 => x"ab",
          8667 => x"a0",
          8668 => x"d4",
          8669 => x"fe",
          8670 => x"59",
          8671 => x"3f",
          8672 => x"53",
          8673 => x"51",
          8674 => x"3f",
          8675 => x"b6",
          8676 => x"e7",
          8677 => x"2e",
          8678 => x"80",
          8679 => x"54",
          8680 => x"53",
          8681 => x"51",
          8682 => x"3f",
          8683 => x"80",
          8684 => x"ff",
          8685 => x"84",
          8686 => x"d2",
          8687 => x"ff",
          8688 => x"86",
          8689 => x"f2",
          8690 => x"1b",
          8691 => x"81",
          8692 => x"52",
          8693 => x"51",
          8694 => x"3f",
          8695 => x"ec",
          8696 => x"9e",
          8697 => x"d4",
          8698 => x"51",
          8699 => x"3f",
          8700 => x"87",
          8701 => x"52",
          8702 => x"9a",
          8703 => x"54",
          8704 => x"7a",
          8705 => x"ff",
          8706 => x"65",
          8707 => x"7a",
          8708 => x"8f",
          8709 => x"80",
          8710 => x"2e",
          8711 => x"9a",
          8712 => x"7a",
          8713 => x"a9",
          8714 => x"84",
          8715 => x"9e",
          8716 => x"0a",
          8717 => x"51",
          8718 => x"ff",
          8719 => x"7d",
          8720 => x"38",
          8721 => x"52",
          8722 => x"9e",
          8723 => x"55",
          8724 => x"62",
          8725 => x"74",
          8726 => x"75",
          8727 => x"7e",
          8728 => x"fe",
          8729 => x"98",
          8730 => x"38",
          8731 => x"82",
          8732 => x"52",
          8733 => x"9e",
          8734 => x"16",
          8735 => x"56",
          8736 => x"38",
          8737 => x"77",
          8738 => x"8d",
          8739 => x"7d",
          8740 => x"38",
          8741 => x"57",
          8742 => x"83",
          8743 => x"76",
          8744 => x"7a",
          8745 => x"ff",
          8746 => x"82",
          8747 => x"81",
          8748 => x"16",
          8749 => x"56",
          8750 => x"38",
          8751 => x"83",
          8752 => x"86",
          8753 => x"ff",
          8754 => x"38",
          8755 => x"82",
          8756 => x"81",
          8757 => x"06",
          8758 => x"fe",
          8759 => x"53",
          8760 => x"51",
          8761 => x"3f",
          8762 => x"52",
          8763 => x"9c",
          8764 => x"be",
          8765 => x"75",
          8766 => x"81",
          8767 => x"0b",
          8768 => x"77",
          8769 => x"75",
          8770 => x"60",
          8771 => x"80",
          8772 => x"75",
          8773 => x"eb",
          8774 => x"85",
          8775 => x"b6",
          8776 => x"2a",
          8777 => x"75",
          8778 => x"82",
          8779 => x"87",
          8780 => x"52",
          8781 => x"51",
          8782 => x"3f",
          8783 => x"ca",
          8784 => x"9c",
          8785 => x"54",
          8786 => x"52",
          8787 => x"98",
          8788 => x"56",
          8789 => x"08",
          8790 => x"53",
          8791 => x"51",
          8792 => x"3f",
          8793 => x"b6",
          8794 => x"38",
          8795 => x"56",
          8796 => x"56",
          8797 => x"b6",
          8798 => x"75",
          8799 => x"0c",
          8800 => x"04",
          8801 => x"7d",
          8802 => x"80",
          8803 => x"05",
          8804 => x"76",
          8805 => x"38",
          8806 => x"11",
          8807 => x"53",
          8808 => x"79",
          8809 => x"3f",
          8810 => x"09",
          8811 => x"38",
          8812 => x"55",
          8813 => x"db",
          8814 => x"70",
          8815 => x"34",
          8816 => x"74",
          8817 => x"81",
          8818 => x"80",
          8819 => x"55",
          8820 => x"76",
          8821 => x"b6",
          8822 => x"3d",
          8823 => x"3d",
          8824 => x"84",
          8825 => x"33",
          8826 => x"8a",
          8827 => x"06",
          8828 => x"52",
          8829 => x"3f",
          8830 => x"56",
          8831 => x"be",
          8832 => x"08",
          8833 => x"05",
          8834 => x"75",
          8835 => x"56",
          8836 => x"a1",
          8837 => x"fc",
          8838 => x"53",
          8839 => x"76",
          8840 => x"dc",
          8841 => x"32",
          8842 => x"72",
          8843 => x"70",
          8844 => x"56",
          8845 => x"18",
          8846 => x"88",
          8847 => x"3d",
          8848 => x"3d",
          8849 => x"11",
          8850 => x"80",
          8851 => x"38",
          8852 => x"05",
          8853 => x"8c",
          8854 => x"08",
          8855 => x"3f",
          8856 => x"08",
          8857 => x"16",
          8858 => x"09",
          8859 => x"38",
          8860 => x"55",
          8861 => x"55",
          8862 => x"98",
          8863 => x"0d",
          8864 => x"0d",
          8865 => x"cc",
          8866 => x"73",
          8867 => x"93",
          8868 => x"0c",
          8869 => x"04",
          8870 => x"02",
          8871 => x"33",
          8872 => x"3d",
          8873 => x"54",
          8874 => x"52",
          8875 => x"ae",
          8876 => x"ff",
          8877 => x"3d",
          8878 => x"00",
          8879 => x"ff",
          8880 => x"ff",
          8881 => x"ff",
          8882 => x"00",
          8883 => x"aa",
          8884 => x"2e",
          8885 => x"35",
          8886 => x"3c",
          8887 => x"43",
          8888 => x"4a",
          8889 => x"51",
          8890 => x"58",
          8891 => x"5f",
          8892 => x"66",
          8893 => x"6d",
          8894 => x"74",
          8895 => x"7a",
          8896 => x"80",
          8897 => x"86",
          8898 => x"8c",
          8899 => x"92",
          8900 => x"98",
          8901 => x"9e",
          8902 => x"a4",
          8903 => x"71",
          8904 => x"77",
          8905 => x"7d",
          8906 => x"83",
          8907 => x"89",
          8908 => x"67",
          8909 => x"67",
          8910 => x"78",
          8911 => x"d0",
          8912 => x"4f",
          8913 => x"3c",
          8914 => x"40",
          8915 => x"a1",
          8916 => x"83",
          8917 => x"19",
          8918 => x"9f",
          8919 => x"22",
          8920 => x"3c",
          8921 => x"78",
          8922 => x"a1",
          8923 => x"40",
          8924 => x"3c",
          8925 => x"3c",
          8926 => x"9f",
          8927 => x"19",
          8928 => x"a1",
          8929 => x"d0",
          8930 => x"31",
          8931 => x"1a",
          8932 => x"1a",
          8933 => x"60",
          8934 => x"1a",
          8935 => x"1a",
          8936 => x"1a",
          8937 => x"1a",
          8938 => x"1a",
          8939 => x"1a",
          8940 => x"1a",
          8941 => x"1d",
          8942 => x"1a",
          8943 => x"48",
          8944 => x"78",
          8945 => x"1a",
          8946 => x"1a",
          8947 => x"1a",
          8948 => x"1a",
          8949 => x"1a",
          8950 => x"1a",
          8951 => x"1a",
          8952 => x"1a",
          8953 => x"1a",
          8954 => x"1a",
          8955 => x"1a",
          8956 => x"1a",
          8957 => x"1a",
          8958 => x"1a",
          8959 => x"1a",
          8960 => x"1a",
          8961 => x"1a",
          8962 => x"1a",
          8963 => x"1a",
          8964 => x"1a",
          8965 => x"1a",
          8966 => x"1a",
          8967 => x"1a",
          8968 => x"1a",
          8969 => x"1a",
          8970 => x"1a",
          8971 => x"1a",
          8972 => x"1a",
          8973 => x"1a",
          8974 => x"1a",
          8975 => x"1a",
          8976 => x"1a",
          8977 => x"1a",
          8978 => x"1a",
          8979 => x"1a",
          8980 => x"1a",
          8981 => x"a8",
          8982 => x"1a",
          8983 => x"1a",
          8984 => x"1a",
          8985 => x"1a",
          8986 => x"16",
          8987 => x"1a",
          8988 => x"1a",
          8989 => x"1a",
          8990 => x"1a",
          8991 => x"1a",
          8992 => x"1a",
          8993 => x"1a",
          8994 => x"1a",
          8995 => x"1a",
          8996 => x"1a",
          8997 => x"d8",
          8998 => x"3f",
          8999 => x"af",
          9000 => x"af",
          9001 => x"af",
          9002 => x"1a",
          9003 => x"3f",
          9004 => x"1a",
          9005 => x"1a",
          9006 => x"98",
          9007 => x"1a",
          9008 => x"1a",
          9009 => x"ec",
          9010 => x"f7",
          9011 => x"1a",
          9012 => x"1a",
          9013 => x"11",
          9014 => x"1a",
          9015 => x"1f",
          9016 => x"1a",
          9017 => x"1a",
          9018 => x"16",
          9019 => x"69",
          9020 => x"00",
          9021 => x"63",
          9022 => x"00",
          9023 => x"69",
          9024 => x"00",
          9025 => x"61",
          9026 => x"00",
          9027 => x"65",
          9028 => x"00",
          9029 => x"65",
          9030 => x"00",
          9031 => x"70",
          9032 => x"00",
          9033 => x"66",
          9034 => x"00",
          9035 => x"6d",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"6c",
          9045 => x"00",
          9046 => x"00",
          9047 => x"74",
          9048 => x"00",
          9049 => x"65",
          9050 => x"00",
          9051 => x"6f",
          9052 => x"00",
          9053 => x"74",
          9054 => x"00",
          9055 => x"73",
          9056 => x"00",
          9057 => x"73",
          9058 => x"00",
          9059 => x"6f",
          9060 => x"00",
          9061 => x"00",
          9062 => x"6b",
          9063 => x"72",
          9064 => x"00",
          9065 => x"65",
          9066 => x"6c",
          9067 => x"72",
          9068 => x"00",
          9069 => x"6b",
          9070 => x"74",
          9071 => x"61",
          9072 => x"00",
          9073 => x"66",
          9074 => x"20",
          9075 => x"6e",
          9076 => x"00",
          9077 => x"70",
          9078 => x"20",
          9079 => x"6e",
          9080 => x"00",
          9081 => x"61",
          9082 => x"20",
          9083 => x"65",
          9084 => x"65",
          9085 => x"00",
          9086 => x"65",
          9087 => x"64",
          9088 => x"65",
          9089 => x"00",
          9090 => x"65",
          9091 => x"72",
          9092 => x"79",
          9093 => x"69",
          9094 => x"2e",
          9095 => x"00",
          9096 => x"65",
          9097 => x"6e",
          9098 => x"20",
          9099 => x"61",
          9100 => x"2e",
          9101 => x"00",
          9102 => x"69",
          9103 => x"72",
          9104 => x"20",
          9105 => x"74",
          9106 => x"65",
          9107 => x"00",
          9108 => x"76",
          9109 => x"75",
          9110 => x"72",
          9111 => x"20",
          9112 => x"61",
          9113 => x"2e",
          9114 => x"00",
          9115 => x"6b",
          9116 => x"74",
          9117 => x"61",
          9118 => x"64",
          9119 => x"00",
          9120 => x"63",
          9121 => x"61",
          9122 => x"6c",
          9123 => x"69",
          9124 => x"79",
          9125 => x"6d",
          9126 => x"75",
          9127 => x"6f",
          9128 => x"69",
          9129 => x"00",
          9130 => x"6d",
          9131 => x"61",
          9132 => x"74",
          9133 => x"00",
          9134 => x"65",
          9135 => x"2c",
          9136 => x"65",
          9137 => x"69",
          9138 => x"63",
          9139 => x"65",
          9140 => x"64",
          9141 => x"00",
          9142 => x"65",
          9143 => x"20",
          9144 => x"6b",
          9145 => x"00",
          9146 => x"75",
          9147 => x"63",
          9148 => x"74",
          9149 => x"6d",
          9150 => x"2e",
          9151 => x"00",
          9152 => x"20",
          9153 => x"79",
          9154 => x"65",
          9155 => x"69",
          9156 => x"2e",
          9157 => x"00",
          9158 => x"61",
          9159 => x"65",
          9160 => x"69",
          9161 => x"72",
          9162 => x"74",
          9163 => x"00",
          9164 => x"63",
          9165 => x"2e",
          9166 => x"00",
          9167 => x"6e",
          9168 => x"20",
          9169 => x"6f",
          9170 => x"00",
          9171 => x"75",
          9172 => x"74",
          9173 => x"25",
          9174 => x"74",
          9175 => x"75",
          9176 => x"74",
          9177 => x"73",
          9178 => x"0a",
          9179 => x"00",
          9180 => x"64",
          9181 => x"00",
          9182 => x"30",
          9183 => x"2c",
          9184 => x"25",
          9185 => x"78",
          9186 => x"3d",
          9187 => x"6c",
          9188 => x"5f",
          9189 => x"3d",
          9190 => x"6c",
          9191 => x"30",
          9192 => x"20",
          9193 => x"6c",
          9194 => x"00",
          9195 => x"6c",
          9196 => x"00",
          9197 => x"00",
          9198 => x"58",
          9199 => x"00",
          9200 => x"20",
          9201 => x"20",
          9202 => x"00",
          9203 => x"58",
          9204 => x"00",
          9205 => x"00",
          9206 => x"00",
          9207 => x"00",
          9208 => x"00",
          9209 => x"20",
          9210 => x"28",
          9211 => x"00",
          9212 => x"30",
          9213 => x"30",
          9214 => x"00",
          9215 => x"30",
          9216 => x"00",
          9217 => x"55",
          9218 => x"65",
          9219 => x"30",
          9220 => x"20",
          9221 => x"25",
          9222 => x"2a",
          9223 => x"00",
          9224 => x"20",
          9225 => x"65",
          9226 => x"70",
          9227 => x"61",
          9228 => x"65",
          9229 => x"00",
          9230 => x"65",
          9231 => x"6e",
          9232 => x"72",
          9233 => x"00",
          9234 => x"20",
          9235 => x"65",
          9236 => x"70",
          9237 => x"00",
          9238 => x"54",
          9239 => x"44",
          9240 => x"74",
          9241 => x"75",
          9242 => x"00",
          9243 => x"54",
          9244 => x"52",
          9245 => x"74",
          9246 => x"75",
          9247 => x"00",
          9248 => x"54",
          9249 => x"58",
          9250 => x"74",
          9251 => x"75",
          9252 => x"00",
          9253 => x"54",
          9254 => x"58",
          9255 => x"74",
          9256 => x"75",
          9257 => x"00",
          9258 => x"54",
          9259 => x"58",
          9260 => x"74",
          9261 => x"75",
          9262 => x"00",
          9263 => x"54",
          9264 => x"58",
          9265 => x"74",
          9266 => x"75",
          9267 => x"00",
          9268 => x"74",
          9269 => x"20",
          9270 => x"74",
          9271 => x"72",
          9272 => x"00",
          9273 => x"62",
          9274 => x"67",
          9275 => x"6d",
          9276 => x"2e",
          9277 => x"00",
          9278 => x"6f",
          9279 => x"63",
          9280 => x"74",
          9281 => x"00",
          9282 => x"2e",
          9283 => x"00",
          9284 => x"00",
          9285 => x"6c",
          9286 => x"74",
          9287 => x"6e",
          9288 => x"61",
          9289 => x"65",
          9290 => x"20",
          9291 => x"64",
          9292 => x"20",
          9293 => x"61",
          9294 => x"69",
          9295 => x"20",
          9296 => x"75",
          9297 => x"79",
          9298 => x"00",
          9299 => x"00",
          9300 => x"61",
          9301 => x"67",
          9302 => x"2e",
          9303 => x"00",
          9304 => x"79",
          9305 => x"2e",
          9306 => x"00",
          9307 => x"70",
          9308 => x"6e",
          9309 => x"2e",
          9310 => x"00",
          9311 => x"6c",
          9312 => x"30",
          9313 => x"2d",
          9314 => x"38",
          9315 => x"25",
          9316 => x"29",
          9317 => x"00",
          9318 => x"70",
          9319 => x"6d",
          9320 => x"00",
          9321 => x"6d",
          9322 => x"74",
          9323 => x"00",
          9324 => x"6c",
          9325 => x"30",
          9326 => x"00",
          9327 => x"00",
          9328 => x"6c",
          9329 => x"30",
          9330 => x"00",
          9331 => x"6c",
          9332 => x"30",
          9333 => x"2d",
          9334 => x"00",
          9335 => x"63",
          9336 => x"6e",
          9337 => x"6f",
          9338 => x"40",
          9339 => x"38",
          9340 => x"2e",
          9341 => x"00",
          9342 => x"6c",
          9343 => x"20",
          9344 => x"65",
          9345 => x"25",
          9346 => x"78",
          9347 => x"2e",
          9348 => x"00",
          9349 => x"6c",
          9350 => x"74",
          9351 => x"65",
          9352 => x"6f",
          9353 => x"28",
          9354 => x"2e",
          9355 => x"00",
          9356 => x"74",
          9357 => x"69",
          9358 => x"61",
          9359 => x"69",
          9360 => x"69",
          9361 => x"2e",
          9362 => x"00",
          9363 => x"64",
          9364 => x"62",
          9365 => x"69",
          9366 => x"2e",
          9367 => x"00",
          9368 => x"00",
          9369 => x"00",
          9370 => x"5c",
          9371 => x"25",
          9372 => x"73",
          9373 => x"00",
          9374 => x"5c",
          9375 => x"25",
          9376 => x"00",
          9377 => x"5c",
          9378 => x"00",
          9379 => x"20",
          9380 => x"6d",
          9381 => x"2e",
          9382 => x"00",
          9383 => x"6e",
          9384 => x"2e",
          9385 => x"00",
          9386 => x"62",
          9387 => x"67",
          9388 => x"74",
          9389 => x"75",
          9390 => x"2e",
          9391 => x"00",
          9392 => x"25",
          9393 => x"64",
          9394 => x"3a",
          9395 => x"25",
          9396 => x"64",
          9397 => x"00",
          9398 => x"20",
          9399 => x"66",
          9400 => x"72",
          9401 => x"6f",
          9402 => x"00",
          9403 => x"72",
          9404 => x"53",
          9405 => x"63",
          9406 => x"69",
          9407 => x"00",
          9408 => x"65",
          9409 => x"65",
          9410 => x"6d",
          9411 => x"6d",
          9412 => x"65",
          9413 => x"00",
          9414 => x"20",
          9415 => x"53",
          9416 => x"4d",
          9417 => x"25",
          9418 => x"3a",
          9419 => x"58",
          9420 => x"00",
          9421 => x"20",
          9422 => x"41",
          9423 => x"20",
          9424 => x"25",
          9425 => x"3a",
          9426 => x"58",
          9427 => x"00",
          9428 => x"20",
          9429 => x"4e",
          9430 => x"41",
          9431 => x"25",
          9432 => x"3a",
          9433 => x"58",
          9434 => x"00",
          9435 => x"20",
          9436 => x"4d",
          9437 => x"20",
          9438 => x"25",
          9439 => x"3a",
          9440 => x"58",
          9441 => x"00",
          9442 => x"20",
          9443 => x"20",
          9444 => x"20",
          9445 => x"25",
          9446 => x"3a",
          9447 => x"58",
          9448 => x"00",
          9449 => x"20",
          9450 => x"43",
          9451 => x"20",
          9452 => x"44",
          9453 => x"63",
          9454 => x"3d",
          9455 => x"64",
          9456 => x"00",
          9457 => x"20",
          9458 => x"45",
          9459 => x"20",
          9460 => x"54",
          9461 => x"72",
          9462 => x"3d",
          9463 => x"64",
          9464 => x"00",
          9465 => x"20",
          9466 => x"52",
          9467 => x"52",
          9468 => x"43",
          9469 => x"6e",
          9470 => x"3d",
          9471 => x"64",
          9472 => x"00",
          9473 => x"20",
          9474 => x"48",
          9475 => x"45",
          9476 => x"53",
          9477 => x"00",
          9478 => x"20",
          9479 => x"49",
          9480 => x"00",
          9481 => x"20",
          9482 => x"54",
          9483 => x"00",
          9484 => x"20",
          9485 => x"00",
          9486 => x"20",
          9487 => x"00",
          9488 => x"72",
          9489 => x"65",
          9490 => x"00",
          9491 => x"20",
          9492 => x"20",
          9493 => x"65",
          9494 => x"65",
          9495 => x"72",
          9496 => x"64",
          9497 => x"73",
          9498 => x"25",
          9499 => x"0a",
          9500 => x"00",
          9501 => x"20",
          9502 => x"20",
          9503 => x"6f",
          9504 => x"53",
          9505 => x"74",
          9506 => x"64",
          9507 => x"73",
          9508 => x"25",
          9509 => x"0a",
          9510 => x"00",
          9511 => x"20",
          9512 => x"63",
          9513 => x"74",
          9514 => x"20",
          9515 => x"72",
          9516 => x"20",
          9517 => x"20",
          9518 => x"25",
          9519 => x"0a",
          9520 => x"00",
          9521 => x"63",
          9522 => x"00",
          9523 => x"20",
          9524 => x"20",
          9525 => x"20",
          9526 => x"20",
          9527 => x"20",
          9528 => x"20",
          9529 => x"20",
          9530 => x"25",
          9531 => x"0a",
          9532 => x"00",
          9533 => x"20",
          9534 => x"74",
          9535 => x"43",
          9536 => x"6b",
          9537 => x"65",
          9538 => x"20",
          9539 => x"20",
          9540 => x"25",
          9541 => x"30",
          9542 => x"48",
          9543 => x"00",
          9544 => x"20",
          9545 => x"41",
          9546 => x"6c",
          9547 => x"20",
          9548 => x"71",
          9549 => x"20",
          9550 => x"20",
          9551 => x"25",
          9552 => x"30",
          9553 => x"48",
          9554 => x"00",
          9555 => x"20",
          9556 => x"68",
          9557 => x"65",
          9558 => x"52",
          9559 => x"43",
          9560 => x"6b",
          9561 => x"65",
          9562 => x"25",
          9563 => x"30",
          9564 => x"48",
          9565 => x"00",
          9566 => x"6c",
          9567 => x"00",
          9568 => x"69",
          9569 => x"00",
          9570 => x"78",
          9571 => x"00",
          9572 => x"00",
          9573 => x"6d",
          9574 => x"00",
          9575 => x"6e",
          9576 => x"00",
          9577 => x"00",
          9578 => x"00",
          9579 => x"02",
          9580 => x"fc",
          9581 => x"00",
          9582 => x"03",
          9583 => x"f8",
          9584 => x"00",
          9585 => x"04",
          9586 => x"f4",
          9587 => x"00",
          9588 => x"05",
          9589 => x"f0",
          9590 => x"00",
          9591 => x"06",
          9592 => x"ec",
          9593 => x"00",
          9594 => x"07",
          9595 => x"e8",
          9596 => x"00",
          9597 => x"01",
          9598 => x"e4",
          9599 => x"00",
          9600 => x"08",
          9601 => x"e0",
          9602 => x"00",
          9603 => x"0b",
          9604 => x"dc",
          9605 => x"00",
          9606 => x"09",
          9607 => x"d8",
          9608 => x"00",
          9609 => x"0a",
          9610 => x"d4",
          9611 => x"00",
          9612 => x"0d",
          9613 => x"d0",
          9614 => x"00",
          9615 => x"0c",
          9616 => x"cc",
          9617 => x"00",
          9618 => x"0e",
          9619 => x"c8",
          9620 => x"00",
          9621 => x"0f",
          9622 => x"c4",
          9623 => x"00",
          9624 => x"0f",
          9625 => x"c0",
          9626 => x"00",
          9627 => x"10",
          9628 => x"bc",
          9629 => x"00",
          9630 => x"11",
          9631 => x"b8",
          9632 => x"00",
          9633 => x"12",
          9634 => x"b4",
          9635 => x"00",
          9636 => x"13",
          9637 => x"b0",
          9638 => x"00",
          9639 => x"14",
          9640 => x"ac",
          9641 => x"00",
          9642 => x"15",
          9643 => x"00",
          9644 => x"00",
          9645 => x"00",
          9646 => x"00",
          9647 => x"7e",
          9648 => x"7e",
          9649 => x"7e",
          9650 => x"00",
          9651 => x"7e",
          9652 => x"7e",
          9653 => x"7e",
          9654 => x"00",
          9655 => x"00",
          9656 => x"00",
          9657 => x"00",
          9658 => x"00",
          9659 => x"00",
          9660 => x"00",
          9661 => x"00",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"74",
          9666 => x"00",
          9667 => x"74",
          9668 => x"00",
          9669 => x"00",
          9670 => x"6c",
          9671 => x"25",
          9672 => x"00",
          9673 => x"6c",
          9674 => x"74",
          9675 => x"65",
          9676 => x"20",
          9677 => x"20",
          9678 => x"74",
          9679 => x"20",
          9680 => x"65",
          9681 => x"20",
          9682 => x"2e",
          9683 => x"00",
          9684 => x"6e",
          9685 => x"6f",
          9686 => x"2f",
          9687 => x"61",
          9688 => x"68",
          9689 => x"6f",
          9690 => x"66",
          9691 => x"2c",
          9692 => x"73",
          9693 => x"69",
          9694 => x"00",
          9695 => x"00",
          9696 => x"2c",
          9697 => x"3d",
          9698 => x"5d",
          9699 => x"00",
          9700 => x"00",
          9701 => x"33",
          9702 => x"00",
          9703 => x"4d",
          9704 => x"53",
          9705 => x"00",
          9706 => x"4e",
          9707 => x"20",
          9708 => x"46",
          9709 => x"32",
          9710 => x"00",
          9711 => x"4e",
          9712 => x"20",
          9713 => x"46",
          9714 => x"20",
          9715 => x"00",
          9716 => x"7c",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"41",
          9721 => x"80",
          9722 => x"49",
          9723 => x"8f",
          9724 => x"4f",
          9725 => x"55",
          9726 => x"9b",
          9727 => x"9f",
          9728 => x"55",
          9729 => x"a7",
          9730 => x"ab",
          9731 => x"af",
          9732 => x"b3",
          9733 => x"b7",
          9734 => x"bb",
          9735 => x"bf",
          9736 => x"c3",
          9737 => x"c7",
          9738 => x"cb",
          9739 => x"cf",
          9740 => x"d3",
          9741 => x"d7",
          9742 => x"db",
          9743 => x"df",
          9744 => x"e3",
          9745 => x"e7",
          9746 => x"eb",
          9747 => x"ef",
          9748 => x"f3",
          9749 => x"f7",
          9750 => x"fb",
          9751 => x"ff",
          9752 => x"3b",
          9753 => x"2f",
          9754 => x"3a",
          9755 => x"7c",
          9756 => x"00",
          9757 => x"04",
          9758 => x"40",
          9759 => x"00",
          9760 => x"00",
          9761 => x"02",
          9762 => x"08",
          9763 => x"20",
          9764 => x"00",
          9765 => x"00",
          9766 => x"ec",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"f4",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"fc",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"04",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"0c",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"14",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"1c",
          9791 => x"00",
          9792 => x"00",
          9793 => x"00",
          9794 => x"24",
          9795 => x"00",
          9796 => x"00",
          9797 => x"00",
          9798 => x"2c",
          9799 => x"00",
          9800 => x"00",
          9801 => x"00",
          9802 => x"34",
          9803 => x"00",
          9804 => x"00",
          9805 => x"00",
          9806 => x"38",
          9807 => x"00",
          9808 => x"00",
          9809 => x"00",
          9810 => x"3c",
          9811 => x"00",
          9812 => x"00",
          9813 => x"00",
          9814 => x"40",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"44",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"48",
          9823 => x"00",
          9824 => x"00",
          9825 => x"00",
          9826 => x"4c",
          9827 => x"00",
          9828 => x"00",
          9829 => x"00",
          9830 => x"50",
          9831 => x"00",
          9832 => x"00",
          9833 => x"00",
          9834 => x"58",
          9835 => x"00",
          9836 => x"00",
          9837 => x"00",
          9838 => x"5c",
          9839 => x"00",
          9840 => x"00",
          9841 => x"00",
          9842 => x"64",
          9843 => x"00",
          9844 => x"00",
          9845 => x"00",
          9846 => x"6c",
          9847 => x"00",
          9848 => x"00",
          9849 => x"00",
          9850 => x"74",
          9851 => x"00",
          9852 => x"00",
          9853 => x"00",
          9854 => x"7c",
          9855 => x"00",
          9856 => x"00",
          9857 => x"00",
          9858 => x"84",
          9859 => x"00",
          9860 => x"00",
          9861 => x"00",
          9862 => x"8c",
          9863 => x"00",
          9864 => x"00",
          9865 => x"00",
          9866 => x"94",
          9867 => x"00",
          9868 => x"00",
          9869 => x"00",
          9870 => x"00",
          9871 => x"00",
          9872 => x"ff",
          9873 => x"00",
          9874 => x"ff",
          9875 => x"00",
          9876 => x"ff",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"ff",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"00",
          9886 => x"00",
          9887 => x"00",
          9888 => x"00",
          9889 => x"01",
          9890 => x"01",
          9891 => x"01",
          9892 => x"00",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"00",
          9898 => x"00",
          9899 => x"00",
          9900 => x"00",
          9901 => x"00",
          9902 => x"00",
          9903 => x"00",
          9904 => x"00",
          9905 => x"00",
          9906 => x"00",
          9907 => x"00",
          9908 => x"00",
          9909 => x"00",
          9910 => x"00",
          9911 => x"00",
          9912 => x"00",
          9913 => x"00",
          9914 => x"00",
          9915 => x"00",
          9916 => x"00",
          9917 => x"04",
          9918 => x"00",
          9919 => x"0c",
          9920 => x"00",
          9921 => x"14",
          9922 => x"00",
          9923 => x"00",
          9924 => x"00",
          9925 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"83",
             1 => x"0b",
             2 => x"b9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c2",
           273 => x"0b",
           274 => x"0b",
           275 => x"e0",
           276 => x"0b",
           277 => x"0b",
           278 => x"80",
           279 => x"0b",
           280 => x"0b",
           281 => x"9e",
           282 => x"0b",
           283 => x"0b",
           284 => x"bd",
           285 => x"0b",
           286 => x"0b",
           287 => x"dd",
           288 => x"0b",
           289 => x"0b",
           290 => x"fd",
           291 => x"0b",
           292 => x"0b",
           293 => x"9d",
           294 => x"0b",
           295 => x"0b",
           296 => x"bd",
           297 => x"0b",
           298 => x"0b",
           299 => x"dd",
           300 => x"0b",
           301 => x"0b",
           302 => x"fd",
           303 => x"0b",
           304 => x"0b",
           305 => x"9d",
           306 => x"0b",
           307 => x"0b",
           308 => x"bd",
           309 => x"0b",
           310 => x"0b",
           311 => x"dd",
           312 => x"0b",
           313 => x"0b",
           314 => x"fd",
           315 => x"0b",
           316 => x"0b",
           317 => x"9d",
           318 => x"0b",
           319 => x"0b",
           320 => x"bd",
           321 => x"0b",
           322 => x"0b",
           323 => x"dd",
           324 => x"0b",
           325 => x"0b",
           326 => x"fd",
           327 => x"0b",
           328 => x"0b",
           329 => x"9d",
           330 => x"0b",
           331 => x"0b",
           332 => x"bd",
           333 => x"0b",
           334 => x"0b",
           335 => x"dd",
           336 => x"0b",
           337 => x"0b",
           338 => x"fd",
           339 => x"0b",
           340 => x"0b",
           341 => x"9d",
           342 => x"0b",
           343 => x"0b",
           344 => x"bd",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"b6",
           386 => x"f4",
           387 => x"b6",
           388 => x"d0",
           389 => x"b6",
           390 => x"b2",
           391 => x"a4",
           392 => x"90",
           393 => x"a4",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"82",
           399 => x"82",
           400 => x"82",
           401 => x"94",
           402 => x"b6",
           403 => x"d0",
           404 => x"b6",
           405 => x"c2",
           406 => x"a4",
           407 => x"90",
           408 => x"a4",
           409 => x"cc",
           410 => x"a4",
           411 => x"90",
           412 => x"a4",
           413 => x"fb",
           414 => x"a4",
           415 => x"90",
           416 => x"a4",
           417 => x"2d",
           418 => x"08",
           419 => x"04",
           420 => x"0c",
           421 => x"82",
           422 => x"82",
           423 => x"82",
           424 => x"97",
           425 => x"b6",
           426 => x"d0",
           427 => x"b6",
           428 => x"f8",
           429 => x"b6",
           430 => x"d0",
           431 => x"b6",
           432 => x"f9",
           433 => x"b6",
           434 => x"d0",
           435 => x"b6",
           436 => x"f0",
           437 => x"b6",
           438 => x"d0",
           439 => x"b6",
           440 => x"f2",
           441 => x"b6",
           442 => x"d0",
           443 => x"b6",
           444 => x"f3",
           445 => x"b6",
           446 => x"d0",
           447 => x"b6",
           448 => x"d8",
           449 => x"b6",
           450 => x"d0",
           451 => x"b6",
           452 => x"e5",
           453 => x"b6",
           454 => x"d0",
           455 => x"b6",
           456 => x"dd",
           457 => x"b6",
           458 => x"d0",
           459 => x"b6",
           460 => x"e0",
           461 => x"b6",
           462 => x"d0",
           463 => x"b6",
           464 => x"ea",
           465 => x"b6",
           466 => x"d0",
           467 => x"b6",
           468 => x"f2",
           469 => x"b6",
           470 => x"d0",
           471 => x"b6",
           472 => x"e3",
           473 => x"b6",
           474 => x"d0",
           475 => x"b6",
           476 => x"ed",
           477 => x"b6",
           478 => x"d0",
           479 => x"b6",
           480 => x"ee",
           481 => x"b6",
           482 => x"d0",
           483 => x"b6",
           484 => x"ee",
           485 => x"b6",
           486 => x"d0",
           487 => x"b6",
           488 => x"f6",
           489 => x"b6",
           490 => x"d0",
           491 => x"b6",
           492 => x"f4",
           493 => x"b6",
           494 => x"d0",
           495 => x"b6",
           496 => x"f9",
           497 => x"b6",
           498 => x"d0",
           499 => x"b6",
           500 => x"ef",
           501 => x"b6",
           502 => x"d0",
           503 => x"b6",
           504 => x"fc",
           505 => x"b6",
           506 => x"d0",
           507 => x"b6",
           508 => x"fd",
           509 => x"b6",
           510 => x"d0",
           511 => x"b6",
           512 => x"e5",
           513 => x"b6",
           514 => x"d0",
           515 => x"b6",
           516 => x"e5",
           517 => x"b6",
           518 => x"d0",
           519 => x"b6",
           520 => x"e6",
           521 => x"b6",
           522 => x"d0",
           523 => x"b6",
           524 => x"f0",
           525 => x"b6",
           526 => x"d0",
           527 => x"b6",
           528 => x"fe",
           529 => x"b6",
           530 => x"d0",
           531 => x"b6",
           532 => x"80",
           533 => x"b6",
           534 => x"d0",
           535 => x"b6",
           536 => x"83",
           537 => x"b6",
           538 => x"d0",
           539 => x"b6",
           540 => x"d7",
           541 => x"b6",
           542 => x"d0",
           543 => x"b6",
           544 => x"86",
           545 => x"b6",
           546 => x"d0",
           547 => x"b6",
           548 => x"95",
           549 => x"b6",
           550 => x"d0",
           551 => x"b6",
           552 => x"93",
           553 => x"b6",
           554 => x"d0",
           555 => x"b6",
           556 => x"a8",
           557 => x"b6",
           558 => x"d0",
           559 => x"b6",
           560 => x"aa",
           561 => x"b6",
           562 => x"d0",
           563 => x"b6",
           564 => x"ac",
           565 => x"b6",
           566 => x"d0",
           567 => x"b6",
           568 => x"f0",
           569 => x"b6",
           570 => x"d0",
           571 => x"b6",
           572 => x"f2",
           573 => x"b6",
           574 => x"d0",
           575 => x"b6",
           576 => x"f5",
           577 => x"b6",
           578 => x"d0",
           579 => x"b6",
           580 => x"d6",
           581 => x"b6",
           582 => x"d0",
           583 => x"b6",
           584 => x"a3",
           585 => x"b6",
           586 => x"d0",
           587 => x"b6",
           588 => x"a3",
           589 => x"b6",
           590 => x"d0",
           591 => x"b6",
           592 => x"a7",
           593 => x"b6",
           594 => x"d0",
           595 => x"b6",
           596 => x"9f",
           597 => x"b6",
           598 => x"d0",
           599 => x"04",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"04",
           609 => x"81",
           610 => x"83",
           611 => x"05",
           612 => x"10",
           613 => x"72",
           614 => x"51",
           615 => x"72",
           616 => x"06",
           617 => x"72",
           618 => x"10",
           619 => x"10",
           620 => x"ed",
           621 => x"53",
           622 => x"b6",
           623 => x"cd",
           624 => x"38",
           625 => x"84",
           626 => x"0b",
           627 => x"bc",
           628 => x"51",
           629 => x"04",
           630 => x"a4",
           631 => x"b6",
           632 => x"3d",
           633 => x"a4",
           634 => x"70",
           635 => x"08",
           636 => x"82",
           637 => x"fc",
           638 => x"82",
           639 => x"88",
           640 => x"82",
           641 => x"52",
           642 => x"3f",
           643 => x"08",
           644 => x"a4",
           645 => x"0c",
           646 => x"08",
           647 => x"70",
           648 => x"0c",
           649 => x"3d",
           650 => x"a4",
           651 => x"b6",
           652 => x"82",
           653 => x"fb",
           654 => x"b6",
           655 => x"05",
           656 => x"33",
           657 => x"70",
           658 => x"51",
           659 => x"8f",
           660 => x"82",
           661 => x"8c",
           662 => x"83",
           663 => x"80",
           664 => x"a4",
           665 => x"0c",
           666 => x"82",
           667 => x"8c",
           668 => x"05",
           669 => x"08",
           670 => x"80",
           671 => x"a4",
           672 => x"0c",
           673 => x"08",
           674 => x"82",
           675 => x"fc",
           676 => x"b6",
           677 => x"05",
           678 => x"80",
           679 => x"0b",
           680 => x"08",
           681 => x"25",
           682 => x"82",
           683 => x"90",
           684 => x"a0",
           685 => x"b6",
           686 => x"82",
           687 => x"f8",
           688 => x"82",
           689 => x"f8",
           690 => x"2e",
           691 => x"8d",
           692 => x"82",
           693 => x"f4",
           694 => x"d2",
           695 => x"a4",
           696 => x"08",
           697 => x"08",
           698 => x"53",
           699 => x"34",
           700 => x"08",
           701 => x"ff",
           702 => x"a4",
           703 => x"0c",
           704 => x"08",
           705 => x"81",
           706 => x"a4",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"80",
           711 => x"b6",
           712 => x"05",
           713 => x"b6",
           714 => x"05",
           715 => x"b6",
           716 => x"05",
           717 => x"98",
           718 => x"0d",
           719 => x"0c",
           720 => x"a4",
           721 => x"b6",
           722 => x"3d",
           723 => x"82",
           724 => x"e5",
           725 => x"b6",
           726 => x"05",
           727 => x"a4",
           728 => x"0c",
           729 => x"82",
           730 => x"e8",
           731 => x"b6",
           732 => x"05",
           733 => x"a4",
           734 => x"0c",
           735 => x"08",
           736 => x"54",
           737 => x"08",
           738 => x"53",
           739 => x"08",
           740 => x"53",
           741 => x"8d",
           742 => x"98",
           743 => x"b6",
           744 => x"05",
           745 => x"a4",
           746 => x"08",
           747 => x"08",
           748 => x"05",
           749 => x"74",
           750 => x"a4",
           751 => x"08",
           752 => x"98",
           753 => x"3d",
           754 => x"a4",
           755 => x"b6",
           756 => x"82",
           757 => x"fb",
           758 => x"b6",
           759 => x"05",
           760 => x"a4",
           761 => x"0c",
           762 => x"08",
           763 => x"54",
           764 => x"08",
           765 => x"53",
           766 => x"08",
           767 => x"52",
           768 => x"82",
           769 => x"70",
           770 => x"08",
           771 => x"82",
           772 => x"f8",
           773 => x"82",
           774 => x"51",
           775 => x"0d",
           776 => x"0c",
           777 => x"a4",
           778 => x"b6",
           779 => x"3d",
           780 => x"82",
           781 => x"e4",
           782 => x"b6",
           783 => x"05",
           784 => x"0b",
           785 => x"82",
           786 => x"88",
           787 => x"11",
           788 => x"2a",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"38",
           793 => x"b6",
           794 => x"05",
           795 => x"39",
           796 => x"08",
           797 => x"53",
           798 => x"72",
           799 => x"08",
           800 => x"72",
           801 => x"53",
           802 => x"95",
           803 => x"b6",
           804 => x"05",
           805 => x"82",
           806 => x"8c",
           807 => x"b6",
           808 => x"05",
           809 => x"06",
           810 => x"80",
           811 => x"38",
           812 => x"08",
           813 => x"53",
           814 => x"81",
           815 => x"b6",
           816 => x"05",
           817 => x"b9",
           818 => x"38",
           819 => x"08",
           820 => x"53",
           821 => x"09",
           822 => x"c5",
           823 => x"a4",
           824 => x"33",
           825 => x"70",
           826 => x"51",
           827 => x"38",
           828 => x"08",
           829 => x"70",
           830 => x"81",
           831 => x"06",
           832 => x"53",
           833 => x"99",
           834 => x"a4",
           835 => x"22",
           836 => x"07",
           837 => x"82",
           838 => x"e4",
           839 => x"d0",
           840 => x"a4",
           841 => x"33",
           842 => x"70",
           843 => x"70",
           844 => x"11",
           845 => x"51",
           846 => x"55",
           847 => x"b6",
           848 => x"05",
           849 => x"a4",
           850 => x"33",
           851 => x"a4",
           852 => x"33",
           853 => x"11",
           854 => x"72",
           855 => x"08",
           856 => x"82",
           857 => x"e8",
           858 => x"98",
           859 => x"2c",
           860 => x"72",
           861 => x"38",
           862 => x"82",
           863 => x"e8",
           864 => x"b6",
           865 => x"05",
           866 => x"2a",
           867 => x"51",
           868 => x"fd",
           869 => x"b6",
           870 => x"05",
           871 => x"2b",
           872 => x"70",
           873 => x"88",
           874 => x"51",
           875 => x"82",
           876 => x"ec",
           877 => x"b8",
           878 => x"a4",
           879 => x"22",
           880 => x"70",
           881 => x"51",
           882 => x"2e",
           883 => x"b6",
           884 => x"05",
           885 => x"2b",
           886 => x"51",
           887 => x"8a",
           888 => x"82",
           889 => x"e8",
           890 => x"b6",
           891 => x"05",
           892 => x"82",
           893 => x"c4",
           894 => x"82",
           895 => x"c4",
           896 => x"d8",
           897 => x"38",
           898 => x"08",
           899 => x"70",
           900 => x"97",
           901 => x"08",
           902 => x"53",
           903 => x"b6",
           904 => x"05",
           905 => x"07",
           906 => x"82",
           907 => x"e4",
           908 => x"b6",
           909 => x"05",
           910 => x"07",
           911 => x"82",
           912 => x"e4",
           913 => x"a8",
           914 => x"a4",
           915 => x"22",
           916 => x"07",
           917 => x"82",
           918 => x"e4",
           919 => x"90",
           920 => x"a4",
           921 => x"22",
           922 => x"07",
           923 => x"82",
           924 => x"e4",
           925 => x"f8",
           926 => x"a4",
           927 => x"22",
           928 => x"51",
           929 => x"b6",
           930 => x"05",
           931 => x"82",
           932 => x"e8",
           933 => x"d8",
           934 => x"a4",
           935 => x"22",
           936 => x"51",
           937 => x"b6",
           938 => x"05",
           939 => x"39",
           940 => x"b6",
           941 => x"05",
           942 => x"a4",
           943 => x"22",
           944 => x"53",
           945 => x"a4",
           946 => x"23",
           947 => x"82",
           948 => x"f8",
           949 => x"a8",
           950 => x"a4",
           951 => x"08",
           952 => x"08",
           953 => x"84",
           954 => x"a4",
           955 => x"0c",
           956 => x"53",
           957 => x"a4",
           958 => x"34",
           959 => x"08",
           960 => x"ff",
           961 => x"72",
           962 => x"08",
           963 => x"8c",
           964 => x"b6",
           965 => x"05",
           966 => x"a4",
           967 => x"08",
           968 => x"b6",
           969 => x"05",
           970 => x"82",
           971 => x"fc",
           972 => x"b6",
           973 => x"05",
           974 => x"2a",
           975 => x"51",
           976 => x"72",
           977 => x"38",
           978 => x"08",
           979 => x"70",
           980 => x"72",
           981 => x"82",
           982 => x"fc",
           983 => x"53",
           984 => x"82",
           985 => x"53",
           986 => x"a4",
           987 => x"23",
           988 => x"b6",
           989 => x"05",
           990 => x"8a",
           991 => x"98",
           992 => x"82",
           993 => x"f4",
           994 => x"b6",
           995 => x"05",
           996 => x"b6",
           997 => x"05",
           998 => x"31",
           999 => x"82",
          1000 => x"ec",
          1001 => x"d8",
          1002 => x"a4",
          1003 => x"08",
          1004 => x"08",
          1005 => x"84",
          1006 => x"a4",
          1007 => x"0c",
          1008 => x"b6",
          1009 => x"05",
          1010 => x"a4",
          1011 => x"22",
          1012 => x"70",
          1013 => x"51",
          1014 => x"80",
          1015 => x"82",
          1016 => x"e8",
          1017 => x"98",
          1018 => x"98",
          1019 => x"b6",
          1020 => x"05",
          1021 => x"a1",
          1022 => x"b6",
          1023 => x"72",
          1024 => x"08",
          1025 => x"99",
          1026 => x"a4",
          1027 => x"08",
          1028 => x"3f",
          1029 => x"08",
          1030 => x"b6",
          1031 => x"05",
          1032 => x"a4",
          1033 => x"22",
          1034 => x"a4",
          1035 => x"22",
          1036 => x"54",
          1037 => x"b6",
          1038 => x"05",
          1039 => x"39",
          1040 => x"08",
          1041 => x"70",
          1042 => x"81",
          1043 => x"53",
          1044 => x"a4",
          1045 => x"a4",
          1046 => x"08",
          1047 => x"08",
          1048 => x"84",
          1049 => x"a4",
          1050 => x"0c",
          1051 => x"b6",
          1052 => x"05",
          1053 => x"39",
          1054 => x"08",
          1055 => x"82",
          1056 => x"90",
          1057 => x"05",
          1058 => x"08",
          1059 => x"70",
          1060 => x"a4",
          1061 => x"0c",
          1062 => x"a4",
          1063 => x"08",
          1064 => x"08",
          1065 => x"82",
          1066 => x"fc",
          1067 => x"25",
          1068 => x"b6",
          1069 => x"05",
          1070 => x"07",
          1071 => x"82",
          1072 => x"e4",
          1073 => x"b6",
          1074 => x"05",
          1075 => x"b6",
          1076 => x"05",
          1077 => x"a4",
          1078 => x"22",
          1079 => x"06",
          1080 => x"82",
          1081 => x"e4",
          1082 => x"af",
          1083 => x"82",
          1084 => x"f4",
          1085 => x"39",
          1086 => x"08",
          1087 => x"70",
          1088 => x"51",
          1089 => x"b6",
          1090 => x"05",
          1091 => x"0b",
          1092 => x"08",
          1093 => x"90",
          1094 => x"a4",
          1095 => x"23",
          1096 => x"08",
          1097 => x"70",
          1098 => x"81",
          1099 => x"53",
          1100 => x"a4",
          1101 => x"a4",
          1102 => x"08",
          1103 => x"08",
          1104 => x"84",
          1105 => x"a4",
          1106 => x"0c",
          1107 => x"b6",
          1108 => x"05",
          1109 => x"39",
          1110 => x"08",
          1111 => x"82",
          1112 => x"90",
          1113 => x"05",
          1114 => x"08",
          1115 => x"70",
          1116 => x"a4",
          1117 => x"0c",
          1118 => x"a4",
          1119 => x"08",
          1120 => x"08",
          1121 => x"82",
          1122 => x"e4",
          1123 => x"cf",
          1124 => x"72",
          1125 => x"08",
          1126 => x"82",
          1127 => x"82",
          1128 => x"f0",
          1129 => x"b6",
          1130 => x"05",
          1131 => x"a4",
          1132 => x"22",
          1133 => x"08",
          1134 => x"71",
          1135 => x"56",
          1136 => x"f3",
          1137 => x"98",
          1138 => x"75",
          1139 => x"a4",
          1140 => x"08",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"33",
          1145 => x"73",
          1146 => x"82",
          1147 => x"f0",
          1148 => x"72",
          1149 => x"b6",
          1150 => x"05",
          1151 => x"df",
          1152 => x"53",
          1153 => x"a4",
          1154 => x"34",
          1155 => x"b6",
          1156 => x"05",
          1157 => x"33",
          1158 => x"53",
          1159 => x"a4",
          1160 => x"34",
          1161 => x"08",
          1162 => x"53",
          1163 => x"08",
          1164 => x"73",
          1165 => x"a4",
          1166 => x"08",
          1167 => x"b6",
          1168 => x"05",
          1169 => x"a4",
          1170 => x"22",
          1171 => x"b6",
          1172 => x"05",
          1173 => x"a2",
          1174 => x"b6",
          1175 => x"82",
          1176 => x"fc",
          1177 => x"82",
          1178 => x"fc",
          1179 => x"2e",
          1180 => x"b2",
          1181 => x"a4",
          1182 => x"08",
          1183 => x"54",
          1184 => x"74",
          1185 => x"51",
          1186 => x"b6",
          1187 => x"05",
          1188 => x"a4",
          1189 => x"22",
          1190 => x"51",
          1191 => x"2e",
          1192 => x"b6",
          1193 => x"05",
          1194 => x"51",
          1195 => x"b6",
          1196 => x"05",
          1197 => x"a4",
          1198 => x"22",
          1199 => x"70",
          1200 => x"51",
          1201 => x"2e",
          1202 => x"82",
          1203 => x"ec",
          1204 => x"90",
          1205 => x"a4",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"90",
          1209 => x"a4",
          1210 => x"0c",
          1211 => x"08",
          1212 => x"51",
          1213 => x"2e",
          1214 => x"95",
          1215 => x"a4",
          1216 => x"08",
          1217 => x"72",
          1218 => x"08",
          1219 => x"93",
          1220 => x"a4",
          1221 => x"08",
          1222 => x"72",
          1223 => x"08",
          1224 => x"82",
          1225 => x"c8",
          1226 => x"b6",
          1227 => x"05",
          1228 => x"a4",
          1229 => x"22",
          1230 => x"70",
          1231 => x"51",
          1232 => x"2e",
          1233 => x"82",
          1234 => x"e8",
          1235 => x"98",
          1236 => x"2c",
          1237 => x"08",
          1238 => x"57",
          1239 => x"72",
          1240 => x"38",
          1241 => x"08",
          1242 => x"70",
          1243 => x"53",
          1244 => x"a4",
          1245 => x"23",
          1246 => x"b6",
          1247 => x"05",
          1248 => x"b6",
          1249 => x"05",
          1250 => x"31",
          1251 => x"82",
          1252 => x"e8",
          1253 => x"b6",
          1254 => x"05",
          1255 => x"2a",
          1256 => x"51",
          1257 => x"80",
          1258 => x"82",
          1259 => x"e8",
          1260 => x"88",
          1261 => x"2b",
          1262 => x"70",
          1263 => x"51",
          1264 => x"72",
          1265 => x"a4",
          1266 => x"22",
          1267 => x"51",
          1268 => x"b6",
          1269 => x"05",
          1270 => x"82",
          1271 => x"fc",
          1272 => x"88",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"51",
          1276 => x"72",
          1277 => x"a4",
          1278 => x"22",
          1279 => x"51",
          1280 => x"b6",
          1281 => x"05",
          1282 => x"a4",
          1283 => x"22",
          1284 => x"06",
          1285 => x"b0",
          1286 => x"a4",
          1287 => x"22",
          1288 => x"54",
          1289 => x"a4",
          1290 => x"23",
          1291 => x"70",
          1292 => x"53",
          1293 => x"90",
          1294 => x"a4",
          1295 => x"08",
          1296 => x"8a",
          1297 => x"39",
          1298 => x"08",
          1299 => x"70",
          1300 => x"81",
          1301 => x"53",
          1302 => x"91",
          1303 => x"a4",
          1304 => x"08",
          1305 => x"8a",
          1306 => x"c7",
          1307 => x"a4",
          1308 => x"22",
          1309 => x"70",
          1310 => x"51",
          1311 => x"2e",
          1312 => x"b6",
          1313 => x"05",
          1314 => x"51",
          1315 => x"a3",
          1316 => x"a4",
          1317 => x"22",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"b6",
          1322 => x"05",
          1323 => x"51",
          1324 => x"82",
          1325 => x"e4",
          1326 => x"86",
          1327 => x"06",
          1328 => x"72",
          1329 => x"38",
          1330 => x"08",
          1331 => x"52",
          1332 => x"df",
          1333 => x"a4",
          1334 => x"22",
          1335 => x"2e",
          1336 => x"94",
          1337 => x"a4",
          1338 => x"08",
          1339 => x"a4",
          1340 => x"33",
          1341 => x"3f",
          1342 => x"08",
          1343 => x"70",
          1344 => x"81",
          1345 => x"53",
          1346 => x"b0",
          1347 => x"a4",
          1348 => x"22",
          1349 => x"54",
          1350 => x"a4",
          1351 => x"23",
          1352 => x"70",
          1353 => x"53",
          1354 => x"90",
          1355 => x"a4",
          1356 => x"08",
          1357 => x"88",
          1358 => x"39",
          1359 => x"08",
          1360 => x"70",
          1361 => x"81",
          1362 => x"53",
          1363 => x"b0",
          1364 => x"a4",
          1365 => x"33",
          1366 => x"54",
          1367 => x"a4",
          1368 => x"34",
          1369 => x"70",
          1370 => x"53",
          1371 => x"90",
          1372 => x"a4",
          1373 => x"08",
          1374 => x"88",
          1375 => x"39",
          1376 => x"08",
          1377 => x"70",
          1378 => x"81",
          1379 => x"53",
          1380 => x"82",
          1381 => x"ec",
          1382 => x"11",
          1383 => x"82",
          1384 => x"ec",
          1385 => x"90",
          1386 => x"2c",
          1387 => x"73",
          1388 => x"82",
          1389 => x"88",
          1390 => x"a0",
          1391 => x"3f",
          1392 => x"b6",
          1393 => x"05",
          1394 => x"80",
          1395 => x"81",
          1396 => x"82",
          1397 => x"88",
          1398 => x"82",
          1399 => x"fc",
          1400 => x"87",
          1401 => x"ee",
          1402 => x"a4",
          1403 => x"33",
          1404 => x"f3",
          1405 => x"06",
          1406 => x"82",
          1407 => x"f4",
          1408 => x"11",
          1409 => x"82",
          1410 => x"f4",
          1411 => x"83",
          1412 => x"53",
          1413 => x"ff",
          1414 => x"38",
          1415 => x"08",
          1416 => x"52",
          1417 => x"08",
          1418 => x"70",
          1419 => x"b6",
          1420 => x"05",
          1421 => x"82",
          1422 => x"fc",
          1423 => x"86",
          1424 => x"b7",
          1425 => x"a4",
          1426 => x"33",
          1427 => x"d3",
          1428 => x"06",
          1429 => x"82",
          1430 => x"f4",
          1431 => x"11",
          1432 => x"82",
          1433 => x"f4",
          1434 => x"83",
          1435 => x"53",
          1436 => x"ff",
          1437 => x"38",
          1438 => x"08",
          1439 => x"52",
          1440 => x"08",
          1441 => x"70",
          1442 => x"86",
          1443 => x"b6",
          1444 => x"05",
          1445 => x"82",
          1446 => x"fc",
          1447 => x"b7",
          1448 => x"a4",
          1449 => x"08",
          1450 => x"2e",
          1451 => x"b6",
          1452 => x"05",
          1453 => x"b6",
          1454 => x"05",
          1455 => x"82",
          1456 => x"f0",
          1457 => x"b6",
          1458 => x"05",
          1459 => x"52",
          1460 => x"3f",
          1461 => x"b6",
          1462 => x"05",
          1463 => x"2a",
          1464 => x"51",
          1465 => x"80",
          1466 => x"38",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"72",
          1470 => x"08",
          1471 => x"73",
          1472 => x"90",
          1473 => x"80",
          1474 => x"38",
          1475 => x"08",
          1476 => x"52",
          1477 => x"9b",
          1478 => x"82",
          1479 => x"88",
          1480 => x"82",
          1481 => x"f8",
          1482 => x"85",
          1483 => x"0b",
          1484 => x"08",
          1485 => x"ea",
          1486 => x"b6",
          1487 => x"05",
          1488 => x"a5",
          1489 => x"06",
          1490 => x"0b",
          1491 => x"08",
          1492 => x"80",
          1493 => x"a4",
          1494 => x"23",
          1495 => x"b6",
          1496 => x"05",
          1497 => x"82",
          1498 => x"f4",
          1499 => x"80",
          1500 => x"a4",
          1501 => x"08",
          1502 => x"a4",
          1503 => x"33",
          1504 => x"3f",
          1505 => x"82",
          1506 => x"88",
          1507 => x"11",
          1508 => x"b6",
          1509 => x"05",
          1510 => x"82",
          1511 => x"e0",
          1512 => x"b6",
          1513 => x"3d",
          1514 => x"a4",
          1515 => x"b6",
          1516 => x"82",
          1517 => x"fd",
          1518 => x"cd",
          1519 => x"82",
          1520 => x"8c",
          1521 => x"82",
          1522 => x"88",
          1523 => x"e4",
          1524 => x"b6",
          1525 => x"82",
          1526 => x"54",
          1527 => x"82",
          1528 => x"04",
          1529 => x"08",
          1530 => x"a4",
          1531 => x"0d",
          1532 => x"b6",
          1533 => x"05",
          1534 => x"ec",
          1535 => x"33",
          1536 => x"70",
          1537 => x"81",
          1538 => x"51",
          1539 => x"80",
          1540 => x"ff",
          1541 => x"a4",
          1542 => x"0c",
          1543 => x"82",
          1544 => x"88",
          1545 => x"72",
          1546 => x"a4",
          1547 => x"08",
          1548 => x"b6",
          1549 => x"05",
          1550 => x"82",
          1551 => x"fc",
          1552 => x"81",
          1553 => x"72",
          1554 => x"38",
          1555 => x"08",
          1556 => x"08",
          1557 => x"a4",
          1558 => x"33",
          1559 => x"08",
          1560 => x"2d",
          1561 => x"08",
          1562 => x"2e",
          1563 => x"ff",
          1564 => x"a4",
          1565 => x"0c",
          1566 => x"82",
          1567 => x"82",
          1568 => x"53",
          1569 => x"90",
          1570 => x"72",
          1571 => x"98",
          1572 => x"80",
          1573 => x"ff",
          1574 => x"a4",
          1575 => x"0c",
          1576 => x"08",
          1577 => x"70",
          1578 => x"08",
          1579 => x"53",
          1580 => x"08",
          1581 => x"82",
          1582 => x"87",
          1583 => x"b6",
          1584 => x"82",
          1585 => x"02",
          1586 => x"0c",
          1587 => x"80",
          1588 => x"a4",
          1589 => x"0c",
          1590 => x"08",
          1591 => x"85",
          1592 => x"81",
          1593 => x"32",
          1594 => x"51",
          1595 => x"53",
          1596 => x"8d",
          1597 => x"82",
          1598 => x"f4",
          1599 => x"f3",
          1600 => x"a4",
          1601 => x"08",
          1602 => x"82",
          1603 => x"88",
          1604 => x"05",
          1605 => x"08",
          1606 => x"53",
          1607 => x"a4",
          1608 => x"34",
          1609 => x"06",
          1610 => x"2e",
          1611 => x"b6",
          1612 => x"05",
          1613 => x"a4",
          1614 => x"08",
          1615 => x"a4",
          1616 => x"33",
          1617 => x"08",
          1618 => x"2d",
          1619 => x"08",
          1620 => x"2e",
          1621 => x"ff",
          1622 => x"a4",
          1623 => x"0c",
          1624 => x"82",
          1625 => x"f8",
          1626 => x"82",
          1627 => x"f4",
          1628 => x"82",
          1629 => x"f4",
          1630 => x"b6",
          1631 => x"3d",
          1632 => x"a4",
          1633 => x"b6",
          1634 => x"82",
          1635 => x"fe",
          1636 => x"cd",
          1637 => x"82",
          1638 => x"88",
          1639 => x"93",
          1640 => x"98",
          1641 => x"b6",
          1642 => x"84",
          1643 => x"b6",
          1644 => x"82",
          1645 => x"02",
          1646 => x"0c",
          1647 => x"82",
          1648 => x"8c",
          1649 => x"11",
          1650 => x"2a",
          1651 => x"70",
          1652 => x"51",
          1653 => x"72",
          1654 => x"38",
          1655 => x"b6",
          1656 => x"05",
          1657 => x"39",
          1658 => x"08",
          1659 => x"85",
          1660 => x"82",
          1661 => x"06",
          1662 => x"53",
          1663 => x"80",
          1664 => x"b6",
          1665 => x"05",
          1666 => x"a4",
          1667 => x"08",
          1668 => x"14",
          1669 => x"08",
          1670 => x"82",
          1671 => x"8c",
          1672 => x"08",
          1673 => x"a4",
          1674 => x"08",
          1675 => x"54",
          1676 => x"73",
          1677 => x"74",
          1678 => x"a4",
          1679 => x"08",
          1680 => x"81",
          1681 => x"0c",
          1682 => x"08",
          1683 => x"70",
          1684 => x"08",
          1685 => x"51",
          1686 => x"39",
          1687 => x"08",
          1688 => x"82",
          1689 => x"8c",
          1690 => x"82",
          1691 => x"88",
          1692 => x"81",
          1693 => x"90",
          1694 => x"54",
          1695 => x"82",
          1696 => x"53",
          1697 => x"82",
          1698 => x"8c",
          1699 => x"11",
          1700 => x"8c",
          1701 => x"b6",
          1702 => x"05",
          1703 => x"b6",
          1704 => x"05",
          1705 => x"8a",
          1706 => x"82",
          1707 => x"fc",
          1708 => x"b6",
          1709 => x"05",
          1710 => x"98",
          1711 => x"0d",
          1712 => x"0c",
          1713 => x"a4",
          1714 => x"b6",
          1715 => x"3d",
          1716 => x"a4",
          1717 => x"08",
          1718 => x"70",
          1719 => x"81",
          1720 => x"51",
          1721 => x"2e",
          1722 => x"0b",
          1723 => x"08",
          1724 => x"83",
          1725 => x"b6",
          1726 => x"05",
          1727 => x"33",
          1728 => x"70",
          1729 => x"51",
          1730 => x"80",
          1731 => x"38",
          1732 => x"08",
          1733 => x"82",
          1734 => x"88",
          1735 => x"53",
          1736 => x"70",
          1737 => x"51",
          1738 => x"14",
          1739 => x"a4",
          1740 => x"08",
          1741 => x"81",
          1742 => x"0c",
          1743 => x"08",
          1744 => x"84",
          1745 => x"82",
          1746 => x"f8",
          1747 => x"51",
          1748 => x"39",
          1749 => x"08",
          1750 => x"85",
          1751 => x"82",
          1752 => x"06",
          1753 => x"52",
          1754 => x"80",
          1755 => x"b6",
          1756 => x"05",
          1757 => x"70",
          1758 => x"a4",
          1759 => x"0c",
          1760 => x"b6",
          1761 => x"05",
          1762 => x"82",
          1763 => x"88",
          1764 => x"b6",
          1765 => x"05",
          1766 => x"85",
          1767 => x"a0",
          1768 => x"71",
          1769 => x"ff",
          1770 => x"a4",
          1771 => x"0c",
          1772 => x"82",
          1773 => x"88",
          1774 => x"08",
          1775 => x"0c",
          1776 => x"39",
          1777 => x"08",
          1778 => x"82",
          1779 => x"88",
          1780 => x"94",
          1781 => x"52",
          1782 => x"b6",
          1783 => x"82",
          1784 => x"fc",
          1785 => x"82",
          1786 => x"fc",
          1787 => x"25",
          1788 => x"82",
          1789 => x"88",
          1790 => x"b6",
          1791 => x"05",
          1792 => x"a4",
          1793 => x"08",
          1794 => x"82",
          1795 => x"f0",
          1796 => x"82",
          1797 => x"fc",
          1798 => x"2e",
          1799 => x"95",
          1800 => x"a4",
          1801 => x"08",
          1802 => x"71",
          1803 => x"08",
          1804 => x"93",
          1805 => x"a4",
          1806 => x"08",
          1807 => x"71",
          1808 => x"08",
          1809 => x"82",
          1810 => x"f4",
          1811 => x"82",
          1812 => x"ec",
          1813 => x"13",
          1814 => x"82",
          1815 => x"f8",
          1816 => x"39",
          1817 => x"08",
          1818 => x"8c",
          1819 => x"05",
          1820 => x"82",
          1821 => x"fc",
          1822 => x"81",
          1823 => x"82",
          1824 => x"f8",
          1825 => x"51",
          1826 => x"a4",
          1827 => x"08",
          1828 => x"0c",
          1829 => x"82",
          1830 => x"04",
          1831 => x"08",
          1832 => x"a4",
          1833 => x"0d",
          1834 => x"08",
          1835 => x"82",
          1836 => x"fc",
          1837 => x"b6",
          1838 => x"05",
          1839 => x"a4",
          1840 => x"0c",
          1841 => x"08",
          1842 => x"80",
          1843 => x"38",
          1844 => x"08",
          1845 => x"82",
          1846 => x"fc",
          1847 => x"81",
          1848 => x"b6",
          1849 => x"05",
          1850 => x"a4",
          1851 => x"08",
          1852 => x"b6",
          1853 => x"05",
          1854 => x"81",
          1855 => x"b6",
          1856 => x"05",
          1857 => x"a4",
          1858 => x"08",
          1859 => x"a4",
          1860 => x"0c",
          1861 => x"08",
          1862 => x"82",
          1863 => x"90",
          1864 => x"82",
          1865 => x"f8",
          1866 => x"b6",
          1867 => x"05",
          1868 => x"82",
          1869 => x"90",
          1870 => x"b6",
          1871 => x"05",
          1872 => x"82",
          1873 => x"90",
          1874 => x"b6",
          1875 => x"05",
          1876 => x"81",
          1877 => x"b6",
          1878 => x"05",
          1879 => x"82",
          1880 => x"fc",
          1881 => x"b6",
          1882 => x"05",
          1883 => x"82",
          1884 => x"f8",
          1885 => x"b6",
          1886 => x"05",
          1887 => x"a4",
          1888 => x"08",
          1889 => x"33",
          1890 => x"ae",
          1891 => x"a4",
          1892 => x"08",
          1893 => x"b6",
          1894 => x"05",
          1895 => x"a4",
          1896 => x"08",
          1897 => x"b6",
          1898 => x"05",
          1899 => x"a4",
          1900 => x"08",
          1901 => x"38",
          1902 => x"08",
          1903 => x"51",
          1904 => x"b6",
          1905 => x"05",
          1906 => x"82",
          1907 => x"f8",
          1908 => x"b6",
          1909 => x"05",
          1910 => x"71",
          1911 => x"b6",
          1912 => x"05",
          1913 => x"82",
          1914 => x"fc",
          1915 => x"ad",
          1916 => x"a4",
          1917 => x"08",
          1918 => x"98",
          1919 => x"3d",
          1920 => x"a4",
          1921 => x"b6",
          1922 => x"82",
          1923 => x"fe",
          1924 => x"b6",
          1925 => x"05",
          1926 => x"a4",
          1927 => x"0c",
          1928 => x"08",
          1929 => x"52",
          1930 => x"b6",
          1931 => x"05",
          1932 => x"82",
          1933 => x"fc",
          1934 => x"81",
          1935 => x"51",
          1936 => x"83",
          1937 => x"82",
          1938 => x"fc",
          1939 => x"05",
          1940 => x"08",
          1941 => x"82",
          1942 => x"fc",
          1943 => x"b6",
          1944 => x"05",
          1945 => x"82",
          1946 => x"51",
          1947 => x"82",
          1948 => x"04",
          1949 => x"08",
          1950 => x"a4",
          1951 => x"0d",
          1952 => x"08",
          1953 => x"82",
          1954 => x"fc",
          1955 => x"b6",
          1956 => x"05",
          1957 => x"33",
          1958 => x"08",
          1959 => x"81",
          1960 => x"a4",
          1961 => x"0c",
          1962 => x"08",
          1963 => x"53",
          1964 => x"34",
          1965 => x"08",
          1966 => x"81",
          1967 => x"a4",
          1968 => x"0c",
          1969 => x"06",
          1970 => x"2e",
          1971 => x"be",
          1972 => x"a4",
          1973 => x"08",
          1974 => x"98",
          1975 => x"3d",
          1976 => x"a4",
          1977 => x"b6",
          1978 => x"82",
          1979 => x"fd",
          1980 => x"b6",
          1981 => x"05",
          1982 => x"a4",
          1983 => x"0c",
          1984 => x"08",
          1985 => x"82",
          1986 => x"f8",
          1987 => x"b6",
          1988 => x"05",
          1989 => x"80",
          1990 => x"b6",
          1991 => x"05",
          1992 => x"82",
          1993 => x"90",
          1994 => x"b6",
          1995 => x"05",
          1996 => x"82",
          1997 => x"90",
          1998 => x"b6",
          1999 => x"05",
          2000 => x"ba",
          2001 => x"a4",
          2002 => x"08",
          2003 => x"82",
          2004 => x"f8",
          2005 => x"05",
          2006 => x"08",
          2007 => x"82",
          2008 => x"fc",
          2009 => x"52",
          2010 => x"82",
          2011 => x"fc",
          2012 => x"05",
          2013 => x"08",
          2014 => x"ff",
          2015 => x"b6",
          2016 => x"05",
          2017 => x"b6",
          2018 => x"85",
          2019 => x"b6",
          2020 => x"82",
          2021 => x"02",
          2022 => x"0c",
          2023 => x"82",
          2024 => x"90",
          2025 => x"2e",
          2026 => x"82",
          2027 => x"8c",
          2028 => x"71",
          2029 => x"a4",
          2030 => x"08",
          2031 => x"b6",
          2032 => x"05",
          2033 => x"a4",
          2034 => x"08",
          2035 => x"81",
          2036 => x"54",
          2037 => x"71",
          2038 => x"80",
          2039 => x"b6",
          2040 => x"05",
          2041 => x"33",
          2042 => x"08",
          2043 => x"81",
          2044 => x"a4",
          2045 => x"0c",
          2046 => x"06",
          2047 => x"8d",
          2048 => x"82",
          2049 => x"fc",
          2050 => x"9b",
          2051 => x"a4",
          2052 => x"08",
          2053 => x"b6",
          2054 => x"05",
          2055 => x"a4",
          2056 => x"08",
          2057 => x"38",
          2058 => x"82",
          2059 => x"90",
          2060 => x"2e",
          2061 => x"82",
          2062 => x"88",
          2063 => x"33",
          2064 => x"8d",
          2065 => x"82",
          2066 => x"fc",
          2067 => x"d7",
          2068 => x"a4",
          2069 => x"08",
          2070 => x"b6",
          2071 => x"05",
          2072 => x"a4",
          2073 => x"08",
          2074 => x"52",
          2075 => x"81",
          2076 => x"a4",
          2077 => x"0c",
          2078 => x"b6",
          2079 => x"05",
          2080 => x"82",
          2081 => x"8c",
          2082 => x"33",
          2083 => x"70",
          2084 => x"08",
          2085 => x"53",
          2086 => x"53",
          2087 => x"0b",
          2088 => x"08",
          2089 => x"82",
          2090 => x"fc",
          2091 => x"b6",
          2092 => x"3d",
          2093 => x"a4",
          2094 => x"b6",
          2095 => x"82",
          2096 => x"fd",
          2097 => x"b6",
          2098 => x"05",
          2099 => x"a4",
          2100 => x"0c",
          2101 => x"08",
          2102 => x"8d",
          2103 => x"82",
          2104 => x"fc",
          2105 => x"ec",
          2106 => x"a4",
          2107 => x"08",
          2108 => x"82",
          2109 => x"f8",
          2110 => x"05",
          2111 => x"08",
          2112 => x"70",
          2113 => x"51",
          2114 => x"2e",
          2115 => x"b6",
          2116 => x"05",
          2117 => x"82",
          2118 => x"8c",
          2119 => x"b6",
          2120 => x"05",
          2121 => x"84",
          2122 => x"39",
          2123 => x"08",
          2124 => x"ff",
          2125 => x"a4",
          2126 => x"0c",
          2127 => x"08",
          2128 => x"82",
          2129 => x"88",
          2130 => x"70",
          2131 => x"08",
          2132 => x"51",
          2133 => x"08",
          2134 => x"82",
          2135 => x"85",
          2136 => x"b6",
          2137 => x"82",
          2138 => x"02",
          2139 => x"0c",
          2140 => x"82",
          2141 => x"88",
          2142 => x"b6",
          2143 => x"05",
          2144 => x"a4",
          2145 => x"08",
          2146 => x"d4",
          2147 => x"a4",
          2148 => x"08",
          2149 => x"b6",
          2150 => x"05",
          2151 => x"a4",
          2152 => x"08",
          2153 => x"b6",
          2154 => x"05",
          2155 => x"a4",
          2156 => x"08",
          2157 => x"38",
          2158 => x"08",
          2159 => x"51",
          2160 => x"a4",
          2161 => x"08",
          2162 => x"71",
          2163 => x"a4",
          2164 => x"08",
          2165 => x"b6",
          2166 => x"05",
          2167 => x"39",
          2168 => x"08",
          2169 => x"70",
          2170 => x"0c",
          2171 => x"0d",
          2172 => x"0c",
          2173 => x"a4",
          2174 => x"b6",
          2175 => x"3d",
          2176 => x"82",
          2177 => x"fc",
          2178 => x"b6",
          2179 => x"05",
          2180 => x"b9",
          2181 => x"a4",
          2182 => x"08",
          2183 => x"a4",
          2184 => x"0c",
          2185 => x"b6",
          2186 => x"05",
          2187 => x"a4",
          2188 => x"08",
          2189 => x"0b",
          2190 => x"08",
          2191 => x"82",
          2192 => x"f4",
          2193 => x"b6",
          2194 => x"05",
          2195 => x"a4",
          2196 => x"08",
          2197 => x"38",
          2198 => x"08",
          2199 => x"30",
          2200 => x"08",
          2201 => x"80",
          2202 => x"a4",
          2203 => x"0c",
          2204 => x"08",
          2205 => x"8a",
          2206 => x"82",
          2207 => x"f0",
          2208 => x"b6",
          2209 => x"05",
          2210 => x"a4",
          2211 => x"0c",
          2212 => x"b6",
          2213 => x"05",
          2214 => x"b6",
          2215 => x"05",
          2216 => x"c5",
          2217 => x"98",
          2218 => x"b6",
          2219 => x"05",
          2220 => x"b6",
          2221 => x"05",
          2222 => x"90",
          2223 => x"a4",
          2224 => x"08",
          2225 => x"a4",
          2226 => x"0c",
          2227 => x"08",
          2228 => x"70",
          2229 => x"0c",
          2230 => x"0d",
          2231 => x"0c",
          2232 => x"a4",
          2233 => x"b6",
          2234 => x"3d",
          2235 => x"82",
          2236 => x"fc",
          2237 => x"b6",
          2238 => x"05",
          2239 => x"99",
          2240 => x"a4",
          2241 => x"08",
          2242 => x"a4",
          2243 => x"0c",
          2244 => x"b6",
          2245 => x"05",
          2246 => x"a4",
          2247 => x"08",
          2248 => x"38",
          2249 => x"08",
          2250 => x"30",
          2251 => x"08",
          2252 => x"81",
          2253 => x"a4",
          2254 => x"08",
          2255 => x"a4",
          2256 => x"08",
          2257 => x"3f",
          2258 => x"08",
          2259 => x"a4",
          2260 => x"0c",
          2261 => x"a4",
          2262 => x"08",
          2263 => x"38",
          2264 => x"08",
          2265 => x"30",
          2266 => x"08",
          2267 => x"82",
          2268 => x"f8",
          2269 => x"82",
          2270 => x"54",
          2271 => x"82",
          2272 => x"04",
          2273 => x"08",
          2274 => x"a4",
          2275 => x"0d",
          2276 => x"b6",
          2277 => x"05",
          2278 => x"b6",
          2279 => x"05",
          2280 => x"c5",
          2281 => x"98",
          2282 => x"b6",
          2283 => x"85",
          2284 => x"b6",
          2285 => x"82",
          2286 => x"02",
          2287 => x"0c",
          2288 => x"81",
          2289 => x"a4",
          2290 => x"08",
          2291 => x"a4",
          2292 => x"08",
          2293 => x"82",
          2294 => x"70",
          2295 => x"0c",
          2296 => x"0d",
          2297 => x"0c",
          2298 => x"a4",
          2299 => x"b6",
          2300 => x"3d",
          2301 => x"82",
          2302 => x"fc",
          2303 => x"0b",
          2304 => x"08",
          2305 => x"82",
          2306 => x"8c",
          2307 => x"b6",
          2308 => x"05",
          2309 => x"38",
          2310 => x"08",
          2311 => x"80",
          2312 => x"80",
          2313 => x"a4",
          2314 => x"08",
          2315 => x"82",
          2316 => x"8c",
          2317 => x"82",
          2318 => x"8c",
          2319 => x"b6",
          2320 => x"05",
          2321 => x"b6",
          2322 => x"05",
          2323 => x"39",
          2324 => x"08",
          2325 => x"80",
          2326 => x"38",
          2327 => x"08",
          2328 => x"82",
          2329 => x"88",
          2330 => x"ad",
          2331 => x"a4",
          2332 => x"08",
          2333 => x"08",
          2334 => x"31",
          2335 => x"08",
          2336 => x"82",
          2337 => x"f8",
          2338 => x"b6",
          2339 => x"05",
          2340 => x"b6",
          2341 => x"05",
          2342 => x"a4",
          2343 => x"08",
          2344 => x"b6",
          2345 => x"05",
          2346 => x"a4",
          2347 => x"08",
          2348 => x"b6",
          2349 => x"05",
          2350 => x"39",
          2351 => x"08",
          2352 => x"80",
          2353 => x"82",
          2354 => x"88",
          2355 => x"82",
          2356 => x"f4",
          2357 => x"91",
          2358 => x"a4",
          2359 => x"08",
          2360 => x"a4",
          2361 => x"0c",
          2362 => x"a4",
          2363 => x"08",
          2364 => x"0c",
          2365 => x"82",
          2366 => x"04",
          2367 => x"08",
          2368 => x"a4",
          2369 => x"0d",
          2370 => x"b6",
          2371 => x"05",
          2372 => x"a4",
          2373 => x"08",
          2374 => x"0c",
          2375 => x"08",
          2376 => x"70",
          2377 => x"72",
          2378 => x"82",
          2379 => x"f8",
          2380 => x"81",
          2381 => x"72",
          2382 => x"81",
          2383 => x"82",
          2384 => x"88",
          2385 => x"08",
          2386 => x"0c",
          2387 => x"82",
          2388 => x"f8",
          2389 => x"72",
          2390 => x"81",
          2391 => x"81",
          2392 => x"a4",
          2393 => x"34",
          2394 => x"08",
          2395 => x"70",
          2396 => x"71",
          2397 => x"51",
          2398 => x"82",
          2399 => x"f8",
          2400 => x"b6",
          2401 => x"05",
          2402 => x"b0",
          2403 => x"06",
          2404 => x"82",
          2405 => x"88",
          2406 => x"08",
          2407 => x"0c",
          2408 => x"53",
          2409 => x"b6",
          2410 => x"05",
          2411 => x"a4",
          2412 => x"33",
          2413 => x"08",
          2414 => x"82",
          2415 => x"e8",
          2416 => x"e2",
          2417 => x"82",
          2418 => x"e8",
          2419 => x"f8",
          2420 => x"80",
          2421 => x"0b",
          2422 => x"08",
          2423 => x"82",
          2424 => x"88",
          2425 => x"08",
          2426 => x"0c",
          2427 => x"53",
          2428 => x"b6",
          2429 => x"05",
          2430 => x"39",
          2431 => x"b6",
          2432 => x"05",
          2433 => x"a4",
          2434 => x"08",
          2435 => x"05",
          2436 => x"08",
          2437 => x"33",
          2438 => x"08",
          2439 => x"80",
          2440 => x"b6",
          2441 => x"05",
          2442 => x"a0",
          2443 => x"81",
          2444 => x"a4",
          2445 => x"0c",
          2446 => x"82",
          2447 => x"f8",
          2448 => x"af",
          2449 => x"38",
          2450 => x"08",
          2451 => x"53",
          2452 => x"83",
          2453 => x"80",
          2454 => x"a4",
          2455 => x"0c",
          2456 => x"88",
          2457 => x"a4",
          2458 => x"34",
          2459 => x"b6",
          2460 => x"05",
          2461 => x"73",
          2462 => x"82",
          2463 => x"f8",
          2464 => x"72",
          2465 => x"38",
          2466 => x"0b",
          2467 => x"08",
          2468 => x"82",
          2469 => x"0b",
          2470 => x"08",
          2471 => x"80",
          2472 => x"a4",
          2473 => x"0c",
          2474 => x"08",
          2475 => x"53",
          2476 => x"81",
          2477 => x"b6",
          2478 => x"05",
          2479 => x"e0",
          2480 => x"38",
          2481 => x"08",
          2482 => x"e0",
          2483 => x"72",
          2484 => x"08",
          2485 => x"82",
          2486 => x"f8",
          2487 => x"11",
          2488 => x"82",
          2489 => x"f8",
          2490 => x"b6",
          2491 => x"05",
          2492 => x"73",
          2493 => x"82",
          2494 => x"f8",
          2495 => x"11",
          2496 => x"82",
          2497 => x"f8",
          2498 => x"b6",
          2499 => x"05",
          2500 => x"89",
          2501 => x"80",
          2502 => x"a4",
          2503 => x"0c",
          2504 => x"82",
          2505 => x"f8",
          2506 => x"b6",
          2507 => x"05",
          2508 => x"72",
          2509 => x"38",
          2510 => x"b6",
          2511 => x"05",
          2512 => x"39",
          2513 => x"08",
          2514 => x"70",
          2515 => x"08",
          2516 => x"29",
          2517 => x"08",
          2518 => x"70",
          2519 => x"a4",
          2520 => x"0c",
          2521 => x"08",
          2522 => x"70",
          2523 => x"71",
          2524 => x"51",
          2525 => x"53",
          2526 => x"b6",
          2527 => x"05",
          2528 => x"39",
          2529 => x"08",
          2530 => x"53",
          2531 => x"90",
          2532 => x"a4",
          2533 => x"08",
          2534 => x"a4",
          2535 => x"0c",
          2536 => x"08",
          2537 => x"82",
          2538 => x"fc",
          2539 => x"0c",
          2540 => x"82",
          2541 => x"ec",
          2542 => x"b6",
          2543 => x"05",
          2544 => x"98",
          2545 => x"0d",
          2546 => x"0c",
          2547 => x"a4",
          2548 => x"b6",
          2549 => x"3d",
          2550 => x"82",
          2551 => x"f0",
          2552 => x"b6",
          2553 => x"05",
          2554 => x"73",
          2555 => x"a4",
          2556 => x"08",
          2557 => x"53",
          2558 => x"72",
          2559 => x"08",
          2560 => x"72",
          2561 => x"53",
          2562 => x"09",
          2563 => x"38",
          2564 => x"08",
          2565 => x"70",
          2566 => x"71",
          2567 => x"39",
          2568 => x"08",
          2569 => x"53",
          2570 => x"09",
          2571 => x"38",
          2572 => x"b6",
          2573 => x"05",
          2574 => x"a4",
          2575 => x"08",
          2576 => x"05",
          2577 => x"08",
          2578 => x"33",
          2579 => x"08",
          2580 => x"82",
          2581 => x"f8",
          2582 => x"72",
          2583 => x"81",
          2584 => x"38",
          2585 => x"08",
          2586 => x"70",
          2587 => x"71",
          2588 => x"51",
          2589 => x"82",
          2590 => x"f8",
          2591 => x"b6",
          2592 => x"05",
          2593 => x"a4",
          2594 => x"0c",
          2595 => x"08",
          2596 => x"80",
          2597 => x"38",
          2598 => x"08",
          2599 => x"80",
          2600 => x"38",
          2601 => x"90",
          2602 => x"a4",
          2603 => x"34",
          2604 => x"08",
          2605 => x"70",
          2606 => x"71",
          2607 => x"51",
          2608 => x"82",
          2609 => x"f8",
          2610 => x"a4",
          2611 => x"82",
          2612 => x"f4",
          2613 => x"b6",
          2614 => x"05",
          2615 => x"81",
          2616 => x"70",
          2617 => x"72",
          2618 => x"a4",
          2619 => x"34",
          2620 => x"82",
          2621 => x"f8",
          2622 => x"72",
          2623 => x"38",
          2624 => x"b6",
          2625 => x"05",
          2626 => x"39",
          2627 => x"08",
          2628 => x"53",
          2629 => x"90",
          2630 => x"a4",
          2631 => x"33",
          2632 => x"26",
          2633 => x"39",
          2634 => x"b6",
          2635 => x"05",
          2636 => x"39",
          2637 => x"b6",
          2638 => x"05",
          2639 => x"82",
          2640 => x"f8",
          2641 => x"af",
          2642 => x"38",
          2643 => x"08",
          2644 => x"53",
          2645 => x"83",
          2646 => x"80",
          2647 => x"a4",
          2648 => x"0c",
          2649 => x"8a",
          2650 => x"a4",
          2651 => x"34",
          2652 => x"b6",
          2653 => x"05",
          2654 => x"a4",
          2655 => x"33",
          2656 => x"27",
          2657 => x"82",
          2658 => x"f8",
          2659 => x"80",
          2660 => x"94",
          2661 => x"a4",
          2662 => x"33",
          2663 => x"53",
          2664 => x"a4",
          2665 => x"34",
          2666 => x"08",
          2667 => x"d0",
          2668 => x"72",
          2669 => x"08",
          2670 => x"82",
          2671 => x"f8",
          2672 => x"90",
          2673 => x"38",
          2674 => x"08",
          2675 => x"f9",
          2676 => x"72",
          2677 => x"08",
          2678 => x"82",
          2679 => x"f8",
          2680 => x"72",
          2681 => x"38",
          2682 => x"b6",
          2683 => x"05",
          2684 => x"39",
          2685 => x"08",
          2686 => x"82",
          2687 => x"f4",
          2688 => x"54",
          2689 => x"8d",
          2690 => x"82",
          2691 => x"ec",
          2692 => x"f7",
          2693 => x"a4",
          2694 => x"33",
          2695 => x"a4",
          2696 => x"08",
          2697 => x"a4",
          2698 => x"33",
          2699 => x"b6",
          2700 => x"05",
          2701 => x"a4",
          2702 => x"08",
          2703 => x"05",
          2704 => x"08",
          2705 => x"55",
          2706 => x"82",
          2707 => x"f8",
          2708 => x"a5",
          2709 => x"a4",
          2710 => x"33",
          2711 => x"2e",
          2712 => x"b6",
          2713 => x"05",
          2714 => x"b6",
          2715 => x"05",
          2716 => x"a4",
          2717 => x"08",
          2718 => x"08",
          2719 => x"71",
          2720 => x"0b",
          2721 => x"08",
          2722 => x"82",
          2723 => x"ec",
          2724 => x"b6",
          2725 => x"3d",
          2726 => x"a4",
          2727 => x"3d",
          2728 => x"08",
          2729 => x"58",
          2730 => x"80",
          2731 => x"39",
          2732 => x"e6",
          2733 => x"b6",
          2734 => x"78",
          2735 => x"33",
          2736 => x"39",
          2737 => x"73",
          2738 => x"81",
          2739 => x"81",
          2740 => x"39",
          2741 => x"90",
          2742 => x"98",
          2743 => x"52",
          2744 => x"3f",
          2745 => x"08",
          2746 => x"75",
          2747 => x"a3",
          2748 => x"98",
          2749 => x"84",
          2750 => x"73",
          2751 => x"b0",
          2752 => x"70",
          2753 => x"58",
          2754 => x"27",
          2755 => x"54",
          2756 => x"98",
          2757 => x"0d",
          2758 => x"0d",
          2759 => x"93",
          2760 => x"38",
          2761 => x"82",
          2762 => x"52",
          2763 => x"82",
          2764 => x"81",
          2765 => x"9b",
          2766 => x"f9",
          2767 => x"b4",
          2768 => x"39",
          2769 => x"51",
          2770 => x"82",
          2771 => x"80",
          2772 => x"9b",
          2773 => x"dd",
          2774 => x"f8",
          2775 => x"39",
          2776 => x"51",
          2777 => x"82",
          2778 => x"80",
          2779 => x"9c",
          2780 => x"c1",
          2781 => x"d0",
          2782 => x"82",
          2783 => x"b5",
          2784 => x"80",
          2785 => x"82",
          2786 => x"a9",
          2787 => x"b8",
          2788 => x"82",
          2789 => x"9d",
          2790 => x"e8",
          2791 => x"82",
          2792 => x"91",
          2793 => x"98",
          2794 => x"82",
          2795 => x"85",
          2796 => x"bc",
          2797 => x"3f",
          2798 => x"04",
          2799 => x"77",
          2800 => x"74",
          2801 => x"8a",
          2802 => x"75",
          2803 => x"51",
          2804 => x"e8",
          2805 => x"ef",
          2806 => x"b6",
          2807 => x"75",
          2808 => x"3f",
          2809 => x"08",
          2810 => x"75",
          2811 => x"cc",
          2812 => x"e5",
          2813 => x"0d",
          2814 => x"0d",
          2815 => x"05",
          2816 => x"33",
          2817 => x"68",
          2818 => x"7a",
          2819 => x"51",
          2820 => x"78",
          2821 => x"ff",
          2822 => x"81",
          2823 => x"07",
          2824 => x"06",
          2825 => x"56",
          2826 => x"38",
          2827 => x"52",
          2828 => x"52",
          2829 => x"e7",
          2830 => x"98",
          2831 => x"b6",
          2832 => x"38",
          2833 => x"08",
          2834 => x"88",
          2835 => x"98",
          2836 => x"3d",
          2837 => x"84",
          2838 => x"52",
          2839 => x"84",
          2840 => x"b6",
          2841 => x"82",
          2842 => x"90",
          2843 => x"74",
          2844 => x"38",
          2845 => x"19",
          2846 => x"39",
          2847 => x"05",
          2848 => x"8c",
          2849 => x"70",
          2850 => x"25",
          2851 => x"9f",
          2852 => x"51",
          2853 => x"74",
          2854 => x"38",
          2855 => x"53",
          2856 => x"88",
          2857 => x"51",
          2858 => x"76",
          2859 => x"b6",
          2860 => x"3d",
          2861 => x"3d",
          2862 => x"84",
          2863 => x"33",
          2864 => x"59",
          2865 => x"52",
          2866 => x"ad",
          2867 => x"98",
          2868 => x"38",
          2869 => x"88",
          2870 => x"2e",
          2871 => x"39",
          2872 => x"57",
          2873 => x"56",
          2874 => x"55",
          2875 => x"08",
          2876 => x"ec",
          2877 => x"cd",
          2878 => x"82",
          2879 => x"ff",
          2880 => x"82",
          2881 => x"62",
          2882 => x"82",
          2883 => x"60",
          2884 => x"79",
          2885 => x"98",
          2886 => x"39",
          2887 => x"82",
          2888 => x"8b",
          2889 => x"f3",
          2890 => x"61",
          2891 => x"05",
          2892 => x"33",
          2893 => x"68",
          2894 => x"5c",
          2895 => x"7a",
          2896 => x"ac",
          2897 => x"91",
          2898 => x"b4",
          2899 => x"89",
          2900 => x"74",
          2901 => x"80",
          2902 => x"2e",
          2903 => x"a0",
          2904 => x"80",
          2905 => x"18",
          2906 => x"27",
          2907 => x"22",
          2908 => x"b8",
          2909 => x"e1",
          2910 => x"82",
          2911 => x"ff",
          2912 => x"82",
          2913 => x"c3",
          2914 => x"53",
          2915 => x"8e",
          2916 => x"52",
          2917 => x"51",
          2918 => x"3f",
          2919 => x"9f",
          2920 => x"b8",
          2921 => x"15",
          2922 => x"74",
          2923 => x"7a",
          2924 => x"72",
          2925 => x"9f",
          2926 => x"b8",
          2927 => x"39",
          2928 => x"51",
          2929 => x"3f",
          2930 => x"82",
          2931 => x"52",
          2932 => x"df",
          2933 => x"39",
          2934 => x"51",
          2935 => x"3f",
          2936 => x"79",
          2937 => x"38",
          2938 => x"33",
          2939 => x"56",
          2940 => x"83",
          2941 => x"80",
          2942 => x"27",
          2943 => x"53",
          2944 => x"70",
          2945 => x"51",
          2946 => x"2e",
          2947 => x"80",
          2948 => x"38",
          2949 => x"08",
          2950 => x"88",
          2951 => x"ec",
          2952 => x"51",
          2953 => x"81",
          2954 => x"b6",
          2955 => x"dc",
          2956 => x"3f",
          2957 => x"1c",
          2958 => x"cb",
          2959 => x"98",
          2960 => x"70",
          2961 => x"57",
          2962 => x"09",
          2963 => x"38",
          2964 => x"82",
          2965 => x"98",
          2966 => x"2c",
          2967 => x"70",
          2968 => x"32",
          2969 => x"72",
          2970 => x"07",
          2971 => x"58",
          2972 => x"57",
          2973 => x"d8",
          2974 => x"2e",
          2975 => x"85",
          2976 => x"8c",
          2977 => x"53",
          2978 => x"fd",
          2979 => x"53",
          2980 => x"98",
          2981 => x"0d",
          2982 => x"0d",
          2983 => x"33",
          2984 => x"53",
          2985 => x"52",
          2986 => x"ad",
          2987 => x"f0",
          2988 => x"a4",
          2989 => x"f0",
          2990 => x"fc",
          2991 => x"f1",
          2992 => x"a0",
          2993 => x"b6",
          2994 => x"80",
          2995 => x"a0",
          2996 => x"3d",
          2997 => x"3d",
          2998 => x"96",
          2999 => x"a5",
          3000 => x"51",
          3001 => x"82",
          3002 => x"99",
          3003 => x"51",
          3004 => x"72",
          3005 => x"81",
          3006 => x"71",
          3007 => x"38",
          3008 => x"f0",
          3009 => x"b8",
          3010 => x"3f",
          3011 => x"e4",
          3012 => x"2a",
          3013 => x"51",
          3014 => x"2e",
          3015 => x"51",
          3016 => x"82",
          3017 => x"98",
          3018 => x"51",
          3019 => x"72",
          3020 => x"81",
          3021 => x"71",
          3022 => x"38",
          3023 => x"b4",
          3024 => x"d8",
          3025 => x"3f",
          3026 => x"a8",
          3027 => x"2a",
          3028 => x"51",
          3029 => x"2e",
          3030 => x"51",
          3031 => x"82",
          3032 => x"98",
          3033 => x"51",
          3034 => x"72",
          3035 => x"81",
          3036 => x"71",
          3037 => x"38",
          3038 => x"f8",
          3039 => x"80",
          3040 => x"3f",
          3041 => x"ec",
          3042 => x"2a",
          3043 => x"51",
          3044 => x"2e",
          3045 => x"51",
          3046 => x"82",
          3047 => x"97",
          3048 => x"51",
          3049 => x"72",
          3050 => x"81",
          3051 => x"71",
          3052 => x"38",
          3053 => x"bc",
          3054 => x"a8",
          3055 => x"3f",
          3056 => x"b0",
          3057 => x"2a",
          3058 => x"51",
          3059 => x"2e",
          3060 => x"51",
          3061 => x"82",
          3062 => x"97",
          3063 => x"51",
          3064 => x"a3",
          3065 => x"3d",
          3066 => x"3d",
          3067 => x"84",
          3068 => x"33",
          3069 => x"56",
          3070 => x"51",
          3071 => x"0b",
          3072 => x"94",
          3073 => x"a9",
          3074 => x"82",
          3075 => x"82",
          3076 => x"80",
          3077 => x"82",
          3078 => x"30",
          3079 => x"98",
          3080 => x"25",
          3081 => x"51",
          3082 => x"0b",
          3083 => x"94",
          3084 => x"82",
          3085 => x"54",
          3086 => x"09",
          3087 => x"38",
          3088 => x"53",
          3089 => x"51",
          3090 => x"3f",
          3091 => x"08",
          3092 => x"38",
          3093 => x"08",
          3094 => x"3f",
          3095 => x"cd",
          3096 => x"84",
          3097 => x"0b",
          3098 => x"b1",
          3099 => x"0b",
          3100 => x"33",
          3101 => x"2e",
          3102 => x"8c",
          3103 => x"88",
          3104 => x"75",
          3105 => x"3f",
          3106 => x"b6",
          3107 => x"3d",
          3108 => x"3d",
          3109 => x"71",
          3110 => x"0c",
          3111 => x"52",
          3112 => x"c6",
          3113 => x"b6",
          3114 => x"ff",
          3115 => x"7d",
          3116 => x"06",
          3117 => x"3d",
          3118 => x"82",
          3119 => x"78",
          3120 => x"3f",
          3121 => x"52",
          3122 => x"51",
          3123 => x"3f",
          3124 => x"08",
          3125 => x"38",
          3126 => x"51",
          3127 => x"81",
          3128 => x"82",
          3129 => x"ff",
          3130 => x"96",
          3131 => x"5a",
          3132 => x"79",
          3133 => x"3f",
          3134 => x"84",
          3135 => x"9e",
          3136 => x"98",
          3137 => x"70",
          3138 => x"59",
          3139 => x"2e",
          3140 => x"78",
          3141 => x"b2",
          3142 => x"2e",
          3143 => x"78",
          3144 => x"38",
          3145 => x"ff",
          3146 => x"bc",
          3147 => x"38",
          3148 => x"78",
          3149 => x"83",
          3150 => x"80",
          3151 => x"cd",
          3152 => x"2e",
          3153 => x"8a",
          3154 => x"80",
          3155 => x"d9",
          3156 => x"f9",
          3157 => x"78",
          3158 => x"88",
          3159 => x"80",
          3160 => x"a1",
          3161 => x"39",
          3162 => x"2e",
          3163 => x"78",
          3164 => x"8b",
          3165 => x"82",
          3166 => x"38",
          3167 => x"78",
          3168 => x"89",
          3169 => x"fe",
          3170 => x"ff",
          3171 => x"ff",
          3172 => x"ec",
          3173 => x"b6",
          3174 => x"2e",
          3175 => x"b4",
          3176 => x"11",
          3177 => x"05",
          3178 => x"3f",
          3179 => x"08",
          3180 => x"af",
          3181 => x"fe",
          3182 => x"ff",
          3183 => x"ec",
          3184 => x"b6",
          3185 => x"38",
          3186 => x"08",
          3187 => x"d0",
          3188 => x"85",
          3189 => x"5c",
          3190 => x"27",
          3191 => x"61",
          3192 => x"70",
          3193 => x"0c",
          3194 => x"f5",
          3195 => x"39",
          3196 => x"80",
          3197 => x"84",
          3198 => x"d1",
          3199 => x"98",
          3200 => x"fd",
          3201 => x"3d",
          3202 => x"53",
          3203 => x"51",
          3204 => x"82",
          3205 => x"80",
          3206 => x"38",
          3207 => x"f8",
          3208 => x"84",
          3209 => x"a5",
          3210 => x"98",
          3211 => x"fd",
          3212 => x"a2",
          3213 => x"af",
          3214 => x"5a",
          3215 => x"81",
          3216 => x"59",
          3217 => x"05",
          3218 => x"34",
          3219 => x"42",
          3220 => x"3d",
          3221 => x"53",
          3222 => x"51",
          3223 => x"82",
          3224 => x"80",
          3225 => x"38",
          3226 => x"fc",
          3227 => x"84",
          3228 => x"d9",
          3229 => x"98",
          3230 => x"fc",
          3231 => x"3d",
          3232 => x"53",
          3233 => x"51",
          3234 => x"82",
          3235 => x"80",
          3236 => x"38",
          3237 => x"51",
          3238 => x"3f",
          3239 => x"63",
          3240 => x"61",
          3241 => x"33",
          3242 => x"78",
          3243 => x"38",
          3244 => x"54",
          3245 => x"79",
          3246 => x"fc",
          3247 => x"99",
          3248 => x"62",
          3249 => x"5a",
          3250 => x"51",
          3251 => x"fc",
          3252 => x"3d",
          3253 => x"53",
          3254 => x"51",
          3255 => x"82",
          3256 => x"80",
          3257 => x"b5",
          3258 => x"78",
          3259 => x"38",
          3260 => x"08",
          3261 => x"39",
          3262 => x"33",
          3263 => x"2e",
          3264 => x"b4",
          3265 => x"bc",
          3266 => x"86",
          3267 => x"80",
          3268 => x"82",
          3269 => x"44",
          3270 => x"b5",
          3271 => x"78",
          3272 => x"38",
          3273 => x"08",
          3274 => x"82",
          3275 => x"59",
          3276 => x"88",
          3277 => x"dc",
          3278 => x"39",
          3279 => x"08",
          3280 => x"44",
          3281 => x"fc",
          3282 => x"84",
          3283 => x"fd",
          3284 => x"98",
          3285 => x"38",
          3286 => x"33",
          3287 => x"2e",
          3288 => x"b4",
          3289 => x"80",
          3290 => x"b5",
          3291 => x"78",
          3292 => x"38",
          3293 => x"08",
          3294 => x"82",
          3295 => x"59",
          3296 => x"88",
          3297 => x"d0",
          3298 => x"39",
          3299 => x"33",
          3300 => x"2e",
          3301 => x"b4",
          3302 => x"99",
          3303 => x"82",
          3304 => x"80",
          3305 => x"82",
          3306 => x"43",
          3307 => x"b4",
          3308 => x"05",
          3309 => x"fe",
          3310 => x"ff",
          3311 => x"e8",
          3312 => x"b6",
          3313 => x"2e",
          3314 => x"62",
          3315 => x"88",
          3316 => x"81",
          3317 => x"32",
          3318 => x"72",
          3319 => x"70",
          3320 => x"51",
          3321 => x"80",
          3322 => x"7a",
          3323 => x"38",
          3324 => x"a3",
          3325 => x"ec",
          3326 => x"63",
          3327 => x"62",
          3328 => x"f2",
          3329 => x"a3",
          3330 => x"f5",
          3331 => x"ff",
          3332 => x"ff",
          3333 => x"e7",
          3334 => x"b6",
          3335 => x"2e",
          3336 => x"b4",
          3337 => x"11",
          3338 => x"05",
          3339 => x"3f",
          3340 => x"08",
          3341 => x"38",
          3342 => x"80",
          3343 => x"79",
          3344 => x"05",
          3345 => x"fe",
          3346 => x"ff",
          3347 => x"e6",
          3348 => x"b6",
          3349 => x"38",
          3350 => x"63",
          3351 => x"52",
          3352 => x"51",
          3353 => x"3f",
          3354 => x"08",
          3355 => x"52",
          3356 => x"ab",
          3357 => x"45",
          3358 => x"78",
          3359 => x"e3",
          3360 => x"27",
          3361 => x"3d",
          3362 => x"53",
          3363 => x"51",
          3364 => x"82",
          3365 => x"80",
          3366 => x"63",
          3367 => x"cb",
          3368 => x"34",
          3369 => x"44",
          3370 => x"82",
          3371 => x"c6",
          3372 => x"a7",
          3373 => x"fe",
          3374 => x"ff",
          3375 => x"e0",
          3376 => x"b6",
          3377 => x"2e",
          3378 => x"b4",
          3379 => x"11",
          3380 => x"05",
          3381 => x"3f",
          3382 => x"08",
          3383 => x"38",
          3384 => x"be",
          3385 => x"70",
          3386 => x"23",
          3387 => x"3d",
          3388 => x"53",
          3389 => x"51",
          3390 => x"82",
          3391 => x"e0",
          3392 => x"39",
          3393 => x"54",
          3394 => x"c0",
          3395 => x"c9",
          3396 => x"e8",
          3397 => x"f8",
          3398 => x"ff",
          3399 => x"79",
          3400 => x"59",
          3401 => x"f7",
          3402 => x"9f",
          3403 => x"60",
          3404 => x"d0",
          3405 => x"fe",
          3406 => x"ff",
          3407 => x"df",
          3408 => x"b6",
          3409 => x"2e",
          3410 => x"59",
          3411 => x"22",
          3412 => x"05",
          3413 => x"41",
          3414 => x"82",
          3415 => x"c5",
          3416 => x"a0",
          3417 => x"fe",
          3418 => x"ff",
          3419 => x"df",
          3420 => x"b6",
          3421 => x"2e",
          3422 => x"b4",
          3423 => x"11",
          3424 => x"05",
          3425 => x"3f",
          3426 => x"08",
          3427 => x"38",
          3428 => x"0c",
          3429 => x"05",
          3430 => x"fe",
          3431 => x"ff",
          3432 => x"de",
          3433 => x"b6",
          3434 => x"38",
          3435 => x"60",
          3436 => x"52",
          3437 => x"51",
          3438 => x"3f",
          3439 => x"08",
          3440 => x"52",
          3441 => x"a8",
          3442 => x"45",
          3443 => x"78",
          3444 => x"8f",
          3445 => x"27",
          3446 => x"3d",
          3447 => x"53",
          3448 => x"51",
          3449 => x"82",
          3450 => x"80",
          3451 => x"60",
          3452 => x"59",
          3453 => x"41",
          3454 => x"82",
          3455 => x"c3",
          3456 => x"ab",
          3457 => x"ff",
          3458 => x"ff",
          3459 => x"e3",
          3460 => x"b6",
          3461 => x"2e",
          3462 => x"63",
          3463 => x"dc",
          3464 => x"b5",
          3465 => x"78",
          3466 => x"ff",
          3467 => x"ff",
          3468 => x"e3",
          3469 => x"b6",
          3470 => x"2e",
          3471 => x"63",
          3472 => x"f8",
          3473 => x"91",
          3474 => x"78",
          3475 => x"98",
          3476 => x"f5",
          3477 => x"b6",
          3478 => x"82",
          3479 => x"ff",
          3480 => x"f4",
          3481 => x"a4",
          3482 => x"f8",
          3483 => x"ca",
          3484 => x"39",
          3485 => x"51",
          3486 => x"80",
          3487 => x"39",
          3488 => x"f4",
          3489 => x"45",
          3490 => x"78",
          3491 => x"d3",
          3492 => x"06",
          3493 => x"2e",
          3494 => x"b4",
          3495 => x"05",
          3496 => x"3f",
          3497 => x"08",
          3498 => x"7a",
          3499 => x"38",
          3500 => x"89",
          3501 => x"2e",
          3502 => x"ca",
          3503 => x"2e",
          3504 => x"c2",
          3505 => x"e0",
          3506 => x"82",
          3507 => x"80",
          3508 => x"e8",
          3509 => x"ff",
          3510 => x"ff",
          3511 => x"b8",
          3512 => x"b4",
          3513 => x"05",
          3514 => x"3f",
          3515 => x"55",
          3516 => x"54",
          3517 => x"a4",
          3518 => x"3d",
          3519 => x"51",
          3520 => x"3f",
          3521 => x"54",
          3522 => x"a5",
          3523 => x"3d",
          3524 => x"51",
          3525 => x"3f",
          3526 => x"58",
          3527 => x"57",
          3528 => x"55",
          3529 => x"d0",
          3530 => x"d0",
          3531 => x"3d",
          3532 => x"51",
          3533 => x"82",
          3534 => x"82",
          3535 => x"09",
          3536 => x"72",
          3537 => x"51",
          3538 => x"80",
          3539 => x"26",
          3540 => x"5a",
          3541 => x"59",
          3542 => x"8d",
          3543 => x"70",
          3544 => x"5c",
          3545 => x"c3",
          3546 => x"32",
          3547 => x"07",
          3548 => x"38",
          3549 => x"09",
          3550 => x"e7",
          3551 => x"8c",
          3552 => x"3f",
          3553 => x"f5",
          3554 => x"0b",
          3555 => x"34",
          3556 => x"8c",
          3557 => x"55",
          3558 => x"52",
          3559 => x"e4",
          3560 => x"98",
          3561 => x"75",
          3562 => x"87",
          3563 => x"73",
          3564 => x"3f",
          3565 => x"98",
          3566 => x"0c",
          3567 => x"9c",
          3568 => x"55",
          3569 => x"52",
          3570 => x"b8",
          3571 => x"98",
          3572 => x"75",
          3573 => x"87",
          3574 => x"73",
          3575 => x"3f",
          3576 => x"98",
          3577 => x"0c",
          3578 => x"0b",
          3579 => x"84",
          3580 => x"83",
          3581 => x"94",
          3582 => x"f6",
          3583 => x"f8",
          3584 => x"02",
          3585 => x"05",
          3586 => x"82",
          3587 => x"87",
          3588 => x"13",
          3589 => x"0c",
          3590 => x"0c",
          3591 => x"3f",
          3592 => x"82",
          3593 => x"ff",
          3594 => x"82",
          3595 => x"ff",
          3596 => x"80",
          3597 => x"92",
          3598 => x"51",
          3599 => x"f0",
          3600 => x"04",
          3601 => x"80",
          3602 => x"71",
          3603 => x"87",
          3604 => x"b6",
          3605 => x"ff",
          3606 => x"ff",
          3607 => x"72",
          3608 => x"38",
          3609 => x"98",
          3610 => x"0d",
          3611 => x"0d",
          3612 => x"54",
          3613 => x"52",
          3614 => x"2e",
          3615 => x"72",
          3616 => x"a0",
          3617 => x"06",
          3618 => x"13",
          3619 => x"72",
          3620 => x"a2",
          3621 => x"06",
          3622 => x"13",
          3623 => x"72",
          3624 => x"2e",
          3625 => x"9f",
          3626 => x"81",
          3627 => x"72",
          3628 => x"70",
          3629 => x"38",
          3630 => x"80",
          3631 => x"73",
          3632 => x"39",
          3633 => x"80",
          3634 => x"54",
          3635 => x"83",
          3636 => x"70",
          3637 => x"38",
          3638 => x"80",
          3639 => x"54",
          3640 => x"09",
          3641 => x"38",
          3642 => x"a2",
          3643 => x"70",
          3644 => x"07",
          3645 => x"70",
          3646 => x"38",
          3647 => x"81",
          3648 => x"71",
          3649 => x"51",
          3650 => x"98",
          3651 => x"0d",
          3652 => x"0d",
          3653 => x"08",
          3654 => x"38",
          3655 => x"05",
          3656 => x"d7",
          3657 => x"b6",
          3658 => x"38",
          3659 => x"39",
          3660 => x"82",
          3661 => x"86",
          3662 => x"fc",
          3663 => x"82",
          3664 => x"05",
          3665 => x"52",
          3666 => x"81",
          3667 => x"13",
          3668 => x"51",
          3669 => x"9e",
          3670 => x"38",
          3671 => x"51",
          3672 => x"97",
          3673 => x"38",
          3674 => x"51",
          3675 => x"bb",
          3676 => x"38",
          3677 => x"51",
          3678 => x"bb",
          3679 => x"38",
          3680 => x"55",
          3681 => x"87",
          3682 => x"d9",
          3683 => x"22",
          3684 => x"73",
          3685 => x"80",
          3686 => x"0b",
          3687 => x"9c",
          3688 => x"87",
          3689 => x"0c",
          3690 => x"87",
          3691 => x"0c",
          3692 => x"87",
          3693 => x"0c",
          3694 => x"87",
          3695 => x"0c",
          3696 => x"87",
          3697 => x"0c",
          3698 => x"87",
          3699 => x"0c",
          3700 => x"98",
          3701 => x"87",
          3702 => x"0c",
          3703 => x"c0",
          3704 => x"80",
          3705 => x"b6",
          3706 => x"3d",
          3707 => x"3d",
          3708 => x"87",
          3709 => x"5d",
          3710 => x"87",
          3711 => x"08",
          3712 => x"23",
          3713 => x"b8",
          3714 => x"82",
          3715 => x"c0",
          3716 => x"5a",
          3717 => x"34",
          3718 => x"b0",
          3719 => x"84",
          3720 => x"c0",
          3721 => x"5a",
          3722 => x"34",
          3723 => x"a8",
          3724 => x"86",
          3725 => x"c0",
          3726 => x"5c",
          3727 => x"23",
          3728 => x"a0",
          3729 => x"8a",
          3730 => x"7d",
          3731 => x"ff",
          3732 => x"7b",
          3733 => x"06",
          3734 => x"33",
          3735 => x"33",
          3736 => x"33",
          3737 => x"33",
          3738 => x"33",
          3739 => x"ff",
          3740 => x"82",
          3741 => x"ff",
          3742 => x"8f",
          3743 => x"fb",
          3744 => x"9f",
          3745 => x"b4",
          3746 => x"81",
          3747 => x"55",
          3748 => x"94",
          3749 => x"80",
          3750 => x"87",
          3751 => x"51",
          3752 => x"96",
          3753 => x"06",
          3754 => x"70",
          3755 => x"38",
          3756 => x"70",
          3757 => x"51",
          3758 => x"72",
          3759 => x"81",
          3760 => x"70",
          3761 => x"38",
          3762 => x"70",
          3763 => x"51",
          3764 => x"38",
          3765 => x"06",
          3766 => x"94",
          3767 => x"80",
          3768 => x"87",
          3769 => x"52",
          3770 => x"74",
          3771 => x"0c",
          3772 => x"04",
          3773 => x"02",
          3774 => x"70",
          3775 => x"2a",
          3776 => x"70",
          3777 => x"34",
          3778 => x"04",
          3779 => x"02",
          3780 => x"58",
          3781 => x"09",
          3782 => x"38",
          3783 => x"51",
          3784 => x"b4",
          3785 => x"81",
          3786 => x"56",
          3787 => x"84",
          3788 => x"2e",
          3789 => x"c0",
          3790 => x"72",
          3791 => x"2a",
          3792 => x"55",
          3793 => x"80",
          3794 => x"73",
          3795 => x"81",
          3796 => x"72",
          3797 => x"81",
          3798 => x"06",
          3799 => x"80",
          3800 => x"73",
          3801 => x"81",
          3802 => x"72",
          3803 => x"75",
          3804 => x"53",
          3805 => x"80",
          3806 => x"2e",
          3807 => x"c0",
          3808 => x"77",
          3809 => x"0b",
          3810 => x"0c",
          3811 => x"04",
          3812 => x"79",
          3813 => x"33",
          3814 => x"06",
          3815 => x"70",
          3816 => x"fc",
          3817 => x"ff",
          3818 => x"82",
          3819 => x"70",
          3820 => x"59",
          3821 => x"87",
          3822 => x"51",
          3823 => x"86",
          3824 => x"94",
          3825 => x"08",
          3826 => x"70",
          3827 => x"54",
          3828 => x"2e",
          3829 => x"91",
          3830 => x"06",
          3831 => x"d7",
          3832 => x"32",
          3833 => x"51",
          3834 => x"2e",
          3835 => x"93",
          3836 => x"06",
          3837 => x"ff",
          3838 => x"81",
          3839 => x"87",
          3840 => x"52",
          3841 => x"86",
          3842 => x"94",
          3843 => x"72",
          3844 => x"74",
          3845 => x"ff",
          3846 => x"57",
          3847 => x"38",
          3848 => x"98",
          3849 => x"0d",
          3850 => x"0d",
          3851 => x"33",
          3852 => x"06",
          3853 => x"c0",
          3854 => x"72",
          3855 => x"38",
          3856 => x"94",
          3857 => x"70",
          3858 => x"81",
          3859 => x"51",
          3860 => x"e2",
          3861 => x"ff",
          3862 => x"c0",
          3863 => x"70",
          3864 => x"38",
          3865 => x"90",
          3866 => x"70",
          3867 => x"82",
          3868 => x"51",
          3869 => x"04",
          3870 => x"82",
          3871 => x"81",
          3872 => x"b6",
          3873 => x"fe",
          3874 => x"b4",
          3875 => x"81",
          3876 => x"53",
          3877 => x"84",
          3878 => x"2e",
          3879 => x"c0",
          3880 => x"71",
          3881 => x"2a",
          3882 => x"51",
          3883 => x"52",
          3884 => x"a0",
          3885 => x"ff",
          3886 => x"c0",
          3887 => x"70",
          3888 => x"38",
          3889 => x"90",
          3890 => x"70",
          3891 => x"98",
          3892 => x"51",
          3893 => x"98",
          3894 => x"0d",
          3895 => x"0d",
          3896 => x"80",
          3897 => x"2a",
          3898 => x"51",
          3899 => x"84",
          3900 => x"c0",
          3901 => x"82",
          3902 => x"87",
          3903 => x"08",
          3904 => x"0c",
          3905 => x"94",
          3906 => x"c4",
          3907 => x"9e",
          3908 => x"b4",
          3909 => x"c0",
          3910 => x"82",
          3911 => x"87",
          3912 => x"08",
          3913 => x"0c",
          3914 => x"ac",
          3915 => x"d4",
          3916 => x"9e",
          3917 => x"b4",
          3918 => x"c0",
          3919 => x"82",
          3920 => x"87",
          3921 => x"08",
          3922 => x"0c",
          3923 => x"bc",
          3924 => x"e4",
          3925 => x"9e",
          3926 => x"b4",
          3927 => x"c0",
          3928 => x"82",
          3929 => x"87",
          3930 => x"08",
          3931 => x"b4",
          3932 => x"c0",
          3933 => x"82",
          3934 => x"87",
          3935 => x"08",
          3936 => x"0c",
          3937 => x"8c",
          3938 => x"fc",
          3939 => x"82",
          3940 => x"80",
          3941 => x"9e",
          3942 => x"84",
          3943 => x"51",
          3944 => x"80",
          3945 => x"81",
          3946 => x"b5",
          3947 => x"0b",
          3948 => x"90",
          3949 => x"80",
          3950 => x"52",
          3951 => x"2e",
          3952 => x"52",
          3953 => x"82",
          3954 => x"87",
          3955 => x"08",
          3956 => x"0a",
          3957 => x"52",
          3958 => x"83",
          3959 => x"71",
          3960 => x"34",
          3961 => x"c0",
          3962 => x"70",
          3963 => x"06",
          3964 => x"70",
          3965 => x"38",
          3966 => x"82",
          3967 => x"80",
          3968 => x"9e",
          3969 => x"a0",
          3970 => x"51",
          3971 => x"80",
          3972 => x"81",
          3973 => x"b5",
          3974 => x"0b",
          3975 => x"90",
          3976 => x"80",
          3977 => x"52",
          3978 => x"2e",
          3979 => x"52",
          3980 => x"86",
          3981 => x"87",
          3982 => x"08",
          3983 => x"80",
          3984 => x"52",
          3985 => x"83",
          3986 => x"71",
          3987 => x"34",
          3988 => x"c0",
          3989 => x"70",
          3990 => x"06",
          3991 => x"70",
          3992 => x"38",
          3993 => x"82",
          3994 => x"80",
          3995 => x"9e",
          3996 => x"81",
          3997 => x"51",
          3998 => x"80",
          3999 => x"81",
          4000 => x"b5",
          4001 => x"0b",
          4002 => x"90",
          4003 => x"c0",
          4004 => x"52",
          4005 => x"2e",
          4006 => x"52",
          4007 => x"8a",
          4008 => x"87",
          4009 => x"08",
          4010 => x"06",
          4011 => x"70",
          4012 => x"38",
          4013 => x"82",
          4014 => x"87",
          4015 => x"08",
          4016 => x"06",
          4017 => x"51",
          4018 => x"82",
          4019 => x"80",
          4020 => x"9e",
          4021 => x"84",
          4022 => x"52",
          4023 => x"2e",
          4024 => x"52",
          4025 => x"8d",
          4026 => x"9e",
          4027 => x"83",
          4028 => x"84",
          4029 => x"51",
          4030 => x"8e",
          4031 => x"87",
          4032 => x"08",
          4033 => x"51",
          4034 => x"80",
          4035 => x"81",
          4036 => x"b5",
          4037 => x"c0",
          4038 => x"70",
          4039 => x"51",
          4040 => x"90",
          4041 => x"0d",
          4042 => x"0d",
          4043 => x"51",
          4044 => x"3f",
          4045 => x"33",
          4046 => x"2e",
          4047 => x"a5",
          4048 => x"95",
          4049 => x"a6",
          4050 => x"b1",
          4051 => x"b5",
          4052 => x"73",
          4053 => x"38",
          4054 => x"08",
          4055 => x"08",
          4056 => x"82",
          4057 => x"ff",
          4058 => x"82",
          4059 => x"54",
          4060 => x"94",
          4061 => x"d4",
          4062 => x"d8",
          4063 => x"52",
          4064 => x"51",
          4065 => x"3f",
          4066 => x"33",
          4067 => x"2e",
          4068 => x"b4",
          4069 => x"b4",
          4070 => x"54",
          4071 => x"d0",
          4072 => x"b5",
          4073 => x"85",
          4074 => x"80",
          4075 => x"82",
          4076 => x"82",
          4077 => x"11",
          4078 => x"a6",
          4079 => x"94",
          4080 => x"b5",
          4081 => x"73",
          4082 => x"38",
          4083 => x"08",
          4084 => x"08",
          4085 => x"82",
          4086 => x"ff",
          4087 => x"82",
          4088 => x"54",
          4089 => x"8e",
          4090 => x"8c",
          4091 => x"a7",
          4092 => x"93",
          4093 => x"b5",
          4094 => x"73",
          4095 => x"38",
          4096 => x"33",
          4097 => x"c4",
          4098 => x"cd",
          4099 => x"8d",
          4100 => x"80",
          4101 => x"82",
          4102 => x"52",
          4103 => x"51",
          4104 => x"3f",
          4105 => x"33",
          4106 => x"2e",
          4107 => x"a8",
          4108 => x"af",
          4109 => x"b5",
          4110 => x"73",
          4111 => x"38",
          4112 => x"51",
          4113 => x"3f",
          4114 => x"33",
          4115 => x"2e",
          4116 => x"a8",
          4117 => x"af",
          4118 => x"b5",
          4119 => x"73",
          4120 => x"38",
          4121 => x"51",
          4122 => x"3f",
          4123 => x"33",
          4124 => x"2e",
          4125 => x"a8",
          4126 => x"ae",
          4127 => x"a8",
          4128 => x"ae",
          4129 => x"b4",
          4130 => x"82",
          4131 => x"ff",
          4132 => x"82",
          4133 => x"52",
          4134 => x"51",
          4135 => x"3f",
          4136 => x"08",
          4137 => x"9c",
          4138 => x"ad",
          4139 => x"c4",
          4140 => x"b0",
          4141 => x"f0",
          4142 => x"a9",
          4143 => x"92",
          4144 => x"b4",
          4145 => x"bd",
          4146 => x"75",
          4147 => x"3f",
          4148 => x"08",
          4149 => x"29",
          4150 => x"54",
          4151 => x"98",
          4152 => x"a9",
          4153 => x"91",
          4154 => x"b5",
          4155 => x"73",
          4156 => x"38",
          4157 => x"08",
          4158 => x"c0",
          4159 => x"c5",
          4160 => x"b6",
          4161 => x"84",
          4162 => x"71",
          4163 => x"82",
          4164 => x"52",
          4165 => x"51",
          4166 => x"3f",
          4167 => x"33",
          4168 => x"2e",
          4169 => x"b4",
          4170 => x"bd",
          4171 => x"75",
          4172 => x"3f",
          4173 => x"08",
          4174 => x"29",
          4175 => x"54",
          4176 => x"98",
          4177 => x"aa",
          4178 => x"91",
          4179 => x"51",
          4180 => x"3f",
          4181 => x"04",
          4182 => x"02",
          4183 => x"ff",
          4184 => x"84",
          4185 => x"71",
          4186 => x"96",
          4187 => x"71",
          4188 => x"aa",
          4189 => x"39",
          4190 => x"51",
          4191 => x"ab",
          4192 => x"39",
          4193 => x"51",
          4194 => x"ab",
          4195 => x"39",
          4196 => x"51",
          4197 => x"3f",
          4198 => x"04",
          4199 => x"0c",
          4200 => x"87",
          4201 => x"0c",
          4202 => x"94",
          4203 => x"96",
          4204 => x"fd",
          4205 => x"98",
          4206 => x"2c",
          4207 => x"70",
          4208 => x"10",
          4209 => x"2b",
          4210 => x"54",
          4211 => x"0b",
          4212 => x"12",
          4213 => x"71",
          4214 => x"38",
          4215 => x"11",
          4216 => x"84",
          4217 => x"33",
          4218 => x"52",
          4219 => x"2e",
          4220 => x"83",
          4221 => x"72",
          4222 => x"0c",
          4223 => x"04",
          4224 => x"79",
          4225 => x"a3",
          4226 => x"33",
          4227 => x"72",
          4228 => x"38",
          4229 => x"08",
          4230 => x"ff",
          4231 => x"82",
          4232 => x"52",
          4233 => x"af",
          4234 => x"cd",
          4235 => x"88",
          4236 => x"ff",
          4237 => x"ff",
          4238 => x"74",
          4239 => x"ff",
          4240 => x"39",
          4241 => x"8f",
          4242 => x"74",
          4243 => x"0d",
          4244 => x"0d",
          4245 => x"05",
          4246 => x"02",
          4247 => x"05",
          4248 => x"f0",
          4249 => x"29",
          4250 => x"05",
          4251 => x"59",
          4252 => x"59",
          4253 => x"86",
          4254 => x"9a",
          4255 => x"b5",
          4256 => x"84",
          4257 => x"98",
          4258 => x"70",
          4259 => x"5a",
          4260 => x"82",
          4261 => x"75",
          4262 => x"f0",
          4263 => x"29",
          4264 => x"05",
          4265 => x"56",
          4266 => x"2e",
          4267 => x"53",
          4268 => x"51",
          4269 => x"3f",
          4270 => x"33",
          4271 => x"74",
          4272 => x"34",
          4273 => x"06",
          4274 => x"27",
          4275 => x"0b",
          4276 => x"34",
          4277 => x"b6",
          4278 => x"ec",
          4279 => x"80",
          4280 => x"82",
          4281 => x"55",
          4282 => x"8c",
          4283 => x"54",
          4284 => x"52",
          4285 => x"da",
          4286 => x"b5",
          4287 => x"8a",
          4288 => x"95",
          4289 => x"ec",
          4290 => x"dd",
          4291 => x"3d",
          4292 => x"3d",
          4293 => x"98",
          4294 => x"72",
          4295 => x"80",
          4296 => x"71",
          4297 => x"3f",
          4298 => x"ff",
          4299 => x"54",
          4300 => x"25",
          4301 => x"0b",
          4302 => x"34",
          4303 => x"08",
          4304 => x"2e",
          4305 => x"51",
          4306 => x"3f",
          4307 => x"08",
          4308 => x"3f",
          4309 => x"b5",
          4310 => x"3d",
          4311 => x"3d",
          4312 => x"80",
          4313 => x"ec",
          4314 => x"e3",
          4315 => x"b6",
          4316 => x"d3",
          4317 => x"ec",
          4318 => x"f8",
          4319 => x"70",
          4320 => x"8c",
          4321 => x"b6",
          4322 => x"2e",
          4323 => x"51",
          4324 => x"3f",
          4325 => x"08",
          4326 => x"82",
          4327 => x"25",
          4328 => x"b6",
          4329 => x"05",
          4330 => x"55",
          4331 => x"75",
          4332 => x"81",
          4333 => x"98",
          4334 => x"8c",
          4335 => x"ff",
          4336 => x"06",
          4337 => x"a6",
          4338 => x"d9",
          4339 => x"3d",
          4340 => x"08",
          4341 => x"70",
          4342 => x"52",
          4343 => x"08",
          4344 => x"bb",
          4345 => x"98",
          4346 => x"38",
          4347 => x"b5",
          4348 => x"55",
          4349 => x"8b",
          4350 => x"56",
          4351 => x"3f",
          4352 => x"08",
          4353 => x"38",
          4354 => x"b3",
          4355 => x"b6",
          4356 => x"18",
          4357 => x"0b",
          4358 => x"08",
          4359 => x"82",
          4360 => x"ff",
          4361 => x"55",
          4362 => x"34",
          4363 => x"30",
          4364 => x"9f",
          4365 => x"55",
          4366 => x"85",
          4367 => x"ac",
          4368 => x"ec",
          4369 => x"08",
          4370 => x"e1",
          4371 => x"b6",
          4372 => x"2e",
          4373 => x"ae",
          4374 => x"8a",
          4375 => x"77",
          4376 => x"06",
          4377 => x"52",
          4378 => x"b4",
          4379 => x"51",
          4380 => x"3f",
          4381 => x"54",
          4382 => x"08",
          4383 => x"58",
          4384 => x"98",
          4385 => x"0d",
          4386 => x"0d",
          4387 => x"5c",
          4388 => x"57",
          4389 => x"73",
          4390 => x"81",
          4391 => x"78",
          4392 => x"56",
          4393 => x"98",
          4394 => x"70",
          4395 => x"33",
          4396 => x"73",
          4397 => x"81",
          4398 => x"75",
          4399 => x"38",
          4400 => x"88",
          4401 => x"f4",
          4402 => x"52",
          4403 => x"b6",
          4404 => x"98",
          4405 => x"52",
          4406 => x"ff",
          4407 => x"82",
          4408 => x"80",
          4409 => x"15",
          4410 => x"81",
          4411 => x"74",
          4412 => x"38",
          4413 => x"e6",
          4414 => x"81",
          4415 => x"3d",
          4416 => x"f8",
          4417 => x"c5",
          4418 => x"98",
          4419 => x"9a",
          4420 => x"53",
          4421 => x"51",
          4422 => x"82",
          4423 => x"81",
          4424 => x"74",
          4425 => x"54",
          4426 => x"14",
          4427 => x"06",
          4428 => x"74",
          4429 => x"38",
          4430 => x"82",
          4431 => x"8c",
          4432 => x"d3",
          4433 => x"3d",
          4434 => x"08",
          4435 => x"59",
          4436 => x"0b",
          4437 => x"82",
          4438 => x"82",
          4439 => x"55",
          4440 => x"cb",
          4441 => x"b5",
          4442 => x"55",
          4443 => x"81",
          4444 => x"2e",
          4445 => x"81",
          4446 => x"55",
          4447 => x"2e",
          4448 => x"a8",
          4449 => x"3f",
          4450 => x"08",
          4451 => x"0c",
          4452 => x"08",
          4453 => x"92",
          4454 => x"76",
          4455 => x"98",
          4456 => x"cc",
          4457 => x"b6",
          4458 => x"2e",
          4459 => x"ae",
          4460 => x"a4",
          4461 => x"f7",
          4462 => x"98",
          4463 => x"b5",
          4464 => x"80",
          4465 => x"3d",
          4466 => x"81",
          4467 => x"82",
          4468 => x"56",
          4469 => x"08",
          4470 => x"81",
          4471 => x"38",
          4472 => x"08",
          4473 => x"9e",
          4474 => x"98",
          4475 => x"0b",
          4476 => x"08",
          4477 => x"82",
          4478 => x"ff",
          4479 => x"55",
          4480 => x"34",
          4481 => x"81",
          4482 => x"75",
          4483 => x"3f",
          4484 => x"81",
          4485 => x"54",
          4486 => x"83",
          4487 => x"74",
          4488 => x"81",
          4489 => x"38",
          4490 => x"82",
          4491 => x"76",
          4492 => x"b5",
          4493 => x"2e",
          4494 => x"d6",
          4495 => x"5d",
          4496 => x"82",
          4497 => x"98",
          4498 => x"2c",
          4499 => x"ff",
          4500 => x"78",
          4501 => x"82",
          4502 => x"70",
          4503 => x"98",
          4504 => x"c0",
          4505 => x"2b",
          4506 => x"71",
          4507 => x"70",
          4508 => x"ab",
          4509 => x"08",
          4510 => x"51",
          4511 => x"59",
          4512 => x"5d",
          4513 => x"73",
          4514 => x"e9",
          4515 => x"27",
          4516 => x"81",
          4517 => x"81",
          4518 => x"70",
          4519 => x"55",
          4520 => x"80",
          4521 => x"53",
          4522 => x"51",
          4523 => x"82",
          4524 => x"81",
          4525 => x"73",
          4526 => x"38",
          4527 => x"c0",
          4528 => x"b1",
          4529 => x"80",
          4530 => x"80",
          4531 => x"98",
          4532 => x"ff",
          4533 => x"55",
          4534 => x"97",
          4535 => x"74",
          4536 => x"f5",
          4537 => x"b6",
          4538 => x"ff",
          4539 => x"cc",
          4540 => x"80",
          4541 => x"2e",
          4542 => x"81",
          4543 => x"82",
          4544 => x"74",
          4545 => x"98",
          4546 => x"c0",
          4547 => x"2b",
          4548 => x"70",
          4549 => x"82",
          4550 => x"a8",
          4551 => x"51",
          4552 => x"58",
          4553 => x"77",
          4554 => x"06",
          4555 => x"82",
          4556 => x"08",
          4557 => x"0b",
          4558 => x"34",
          4559 => x"cd",
          4560 => x"39",
          4561 => x"c4",
          4562 => x"cd",
          4563 => x"af",
          4564 => x"7d",
          4565 => x"73",
          4566 => x"e1",
          4567 => x"29",
          4568 => x"05",
          4569 => x"04",
          4570 => x"33",
          4571 => x"2e",
          4572 => x"82",
          4573 => x"55",
          4574 => x"ab",
          4575 => x"2b",
          4576 => x"51",
          4577 => x"24",
          4578 => x"1a",
          4579 => x"81",
          4580 => x"81",
          4581 => x"81",
          4582 => x"70",
          4583 => x"cd",
          4584 => x"51",
          4585 => x"82",
          4586 => x"81",
          4587 => x"74",
          4588 => x"34",
          4589 => x"ae",
          4590 => x"34",
          4591 => x"33",
          4592 => x"25",
          4593 => x"14",
          4594 => x"cd",
          4595 => x"cd",
          4596 => x"81",
          4597 => x"81",
          4598 => x"70",
          4599 => x"cd",
          4600 => x"51",
          4601 => x"77",
          4602 => x"82",
          4603 => x"52",
          4604 => x"33",
          4605 => x"a3",
          4606 => x"81",
          4607 => x"81",
          4608 => x"70",
          4609 => x"cd",
          4610 => x"51",
          4611 => x"24",
          4612 => x"cd",
          4613 => x"98",
          4614 => x"2c",
          4615 => x"33",
          4616 => x"56",
          4617 => x"fc",
          4618 => x"cd",
          4619 => x"88",
          4620 => x"ff",
          4621 => x"80",
          4622 => x"80",
          4623 => x"98",
          4624 => x"c8",
          4625 => x"55",
          4626 => x"de",
          4627 => x"39",
          4628 => x"80",
          4629 => x"34",
          4630 => x"53",
          4631 => x"9e",
          4632 => x"9c",
          4633 => x"39",
          4634 => x"33",
          4635 => x"06",
          4636 => x"80",
          4637 => x"38",
          4638 => x"33",
          4639 => x"73",
          4640 => x"34",
          4641 => x"73",
          4642 => x"34",
          4643 => x"08",
          4644 => x"ff",
          4645 => x"82",
          4646 => x"70",
          4647 => x"98",
          4648 => x"c8",
          4649 => x"56",
          4650 => x"25",
          4651 => x"1a",
          4652 => x"33",
          4653 => x"cd",
          4654 => x"73",
          4655 => x"a1",
          4656 => x"81",
          4657 => x"81",
          4658 => x"70",
          4659 => x"cd",
          4660 => x"51",
          4661 => x"24",
          4662 => x"cd",
          4663 => x"a0",
          4664 => x"cf",
          4665 => x"cc",
          4666 => x"2b",
          4667 => x"82",
          4668 => x"57",
          4669 => x"74",
          4670 => x"c1",
          4671 => x"ec",
          4672 => x"51",
          4673 => x"3f",
          4674 => x"0a",
          4675 => x"0a",
          4676 => x"2c",
          4677 => x"33",
          4678 => x"75",
          4679 => x"38",
          4680 => x"82",
          4681 => x"7a",
          4682 => x"74",
          4683 => x"ec",
          4684 => x"51",
          4685 => x"3f",
          4686 => x"52",
          4687 => x"c9",
          4688 => x"98",
          4689 => x"06",
          4690 => x"38",
          4691 => x"33",
          4692 => x"2e",
          4693 => x"53",
          4694 => x"51",
          4695 => x"84",
          4696 => x"34",
          4697 => x"cd",
          4698 => x"0b",
          4699 => x"34",
          4700 => x"98",
          4701 => x"0d",
          4702 => x"cc",
          4703 => x"80",
          4704 => x"38",
          4705 => x"08",
          4706 => x"ff",
          4707 => x"82",
          4708 => x"ff",
          4709 => x"82",
          4710 => x"73",
          4711 => x"54",
          4712 => x"cd",
          4713 => x"cd",
          4714 => x"55",
          4715 => x"f9",
          4716 => x"14",
          4717 => x"cd",
          4718 => x"98",
          4719 => x"2c",
          4720 => x"06",
          4721 => x"74",
          4722 => x"38",
          4723 => x"81",
          4724 => x"34",
          4725 => x"08",
          4726 => x"51",
          4727 => x"3f",
          4728 => x"0a",
          4729 => x"0a",
          4730 => x"2c",
          4731 => x"33",
          4732 => x"75",
          4733 => x"38",
          4734 => x"08",
          4735 => x"ff",
          4736 => x"82",
          4737 => x"70",
          4738 => x"98",
          4739 => x"c8",
          4740 => x"56",
          4741 => x"24",
          4742 => x"82",
          4743 => x"52",
          4744 => x"9f",
          4745 => x"81",
          4746 => x"81",
          4747 => x"70",
          4748 => x"cd",
          4749 => x"51",
          4750 => x"25",
          4751 => x"fd",
          4752 => x"cc",
          4753 => x"ff",
          4754 => x"c8",
          4755 => x"54",
          4756 => x"f7",
          4757 => x"cd",
          4758 => x"81",
          4759 => x"82",
          4760 => x"74",
          4761 => x"52",
          4762 => x"c7",
          4763 => x"cc",
          4764 => x"ff",
          4765 => x"c8",
          4766 => x"54",
          4767 => x"d6",
          4768 => x"39",
          4769 => x"53",
          4770 => x"9e",
          4771 => x"f0",
          4772 => x"82",
          4773 => x"80",
          4774 => x"c8",
          4775 => x"39",
          4776 => x"82",
          4777 => x"55",
          4778 => x"a6",
          4779 => x"ff",
          4780 => x"82",
          4781 => x"82",
          4782 => x"82",
          4783 => x"81",
          4784 => x"05",
          4785 => x"79",
          4786 => x"9a",
          4787 => x"81",
          4788 => x"84",
          4789 => x"98",
          4790 => x"08",
          4791 => x"80",
          4792 => x"74",
          4793 => x"9e",
          4794 => x"98",
          4795 => x"c8",
          4796 => x"98",
          4797 => x"06",
          4798 => x"74",
          4799 => x"ff",
          4800 => x"ff",
          4801 => x"fa",
          4802 => x"55",
          4803 => x"f6",
          4804 => x"51",
          4805 => x"3f",
          4806 => x"93",
          4807 => x"06",
          4808 => x"b5",
          4809 => x"74",
          4810 => x"38",
          4811 => x"a5",
          4812 => x"b6",
          4813 => x"cd",
          4814 => x"b6",
          4815 => x"ff",
          4816 => x"53",
          4817 => x"51",
          4818 => x"3f",
          4819 => x"7a",
          4820 => x"b5",
          4821 => x"08",
          4822 => x"80",
          4823 => x"74",
          4824 => x"a2",
          4825 => x"98",
          4826 => x"c8",
          4827 => x"98",
          4828 => x"06",
          4829 => x"74",
          4830 => x"ff",
          4831 => x"81",
          4832 => x"81",
          4833 => x"89",
          4834 => x"cd",
          4835 => x"7a",
          4836 => x"cc",
          4837 => x"c8",
          4838 => x"51",
          4839 => x"f5",
          4840 => x"cd",
          4841 => x"81",
          4842 => x"cd",
          4843 => x"56",
          4844 => x"27",
          4845 => x"82",
          4846 => x"52",
          4847 => x"73",
          4848 => x"34",
          4849 => x"33",
          4850 => x"9b",
          4851 => x"ed",
          4852 => x"cc",
          4853 => x"80",
          4854 => x"38",
          4855 => x"08",
          4856 => x"ff",
          4857 => x"82",
          4858 => x"ff",
          4859 => x"82",
          4860 => x"f4",
          4861 => x"3d",
          4862 => x"f4",
          4863 => x"90",
          4864 => x"0b",
          4865 => x"23",
          4866 => x"80",
          4867 => x"f4",
          4868 => x"d3",
          4869 => x"90",
          4870 => x"58",
          4871 => x"81",
          4872 => x"15",
          4873 => x"90",
          4874 => x"84",
          4875 => x"85",
          4876 => x"b6",
          4877 => x"77",
          4878 => x"76",
          4879 => x"82",
          4880 => x"82",
          4881 => x"ff",
          4882 => x"80",
          4883 => x"ff",
          4884 => x"88",
          4885 => x"55",
          4886 => x"17",
          4887 => x"17",
          4888 => x"8c",
          4889 => x"29",
          4890 => x"08",
          4891 => x"51",
          4892 => x"82",
          4893 => x"83",
          4894 => x"3d",
          4895 => x"3d",
          4896 => x"81",
          4897 => x"27",
          4898 => x"12",
          4899 => x"11",
          4900 => x"ff",
          4901 => x"51",
          4902 => x"98",
          4903 => x"0d",
          4904 => x"0d",
          4905 => x"22",
          4906 => x"aa",
          4907 => x"05",
          4908 => x"08",
          4909 => x"71",
          4910 => x"2b",
          4911 => x"33",
          4912 => x"71",
          4913 => x"02",
          4914 => x"05",
          4915 => x"ff",
          4916 => x"70",
          4917 => x"51",
          4918 => x"5b",
          4919 => x"54",
          4920 => x"34",
          4921 => x"34",
          4922 => x"08",
          4923 => x"2a",
          4924 => x"82",
          4925 => x"83",
          4926 => x"b6",
          4927 => x"17",
          4928 => x"12",
          4929 => x"2b",
          4930 => x"2b",
          4931 => x"06",
          4932 => x"52",
          4933 => x"83",
          4934 => x"70",
          4935 => x"54",
          4936 => x"12",
          4937 => x"ff",
          4938 => x"83",
          4939 => x"b6",
          4940 => x"56",
          4941 => x"72",
          4942 => x"89",
          4943 => x"fb",
          4944 => x"b6",
          4945 => x"84",
          4946 => x"22",
          4947 => x"72",
          4948 => x"33",
          4949 => x"71",
          4950 => x"83",
          4951 => x"5b",
          4952 => x"52",
          4953 => x"12",
          4954 => x"33",
          4955 => x"07",
          4956 => x"54",
          4957 => x"70",
          4958 => x"73",
          4959 => x"82",
          4960 => x"70",
          4961 => x"33",
          4962 => x"71",
          4963 => x"83",
          4964 => x"59",
          4965 => x"05",
          4966 => x"87",
          4967 => x"88",
          4968 => x"88",
          4969 => x"56",
          4970 => x"13",
          4971 => x"13",
          4972 => x"90",
          4973 => x"33",
          4974 => x"71",
          4975 => x"70",
          4976 => x"06",
          4977 => x"53",
          4978 => x"53",
          4979 => x"70",
          4980 => x"87",
          4981 => x"fa",
          4982 => x"a2",
          4983 => x"b6",
          4984 => x"83",
          4985 => x"70",
          4986 => x"33",
          4987 => x"07",
          4988 => x"15",
          4989 => x"12",
          4990 => x"2b",
          4991 => x"07",
          4992 => x"55",
          4993 => x"57",
          4994 => x"80",
          4995 => x"38",
          4996 => x"ab",
          4997 => x"90",
          4998 => x"70",
          4999 => x"33",
          5000 => x"71",
          5001 => x"74",
          5002 => x"81",
          5003 => x"88",
          5004 => x"83",
          5005 => x"f8",
          5006 => x"54",
          5007 => x"58",
          5008 => x"74",
          5009 => x"52",
          5010 => x"34",
          5011 => x"34",
          5012 => x"08",
          5013 => x"33",
          5014 => x"71",
          5015 => x"83",
          5016 => x"59",
          5017 => x"05",
          5018 => x"12",
          5019 => x"2b",
          5020 => x"ff",
          5021 => x"88",
          5022 => x"52",
          5023 => x"74",
          5024 => x"15",
          5025 => x"0d",
          5026 => x"0d",
          5027 => x"08",
          5028 => x"9e",
          5029 => x"83",
          5030 => x"82",
          5031 => x"12",
          5032 => x"2b",
          5033 => x"07",
          5034 => x"52",
          5035 => x"05",
          5036 => x"13",
          5037 => x"2b",
          5038 => x"05",
          5039 => x"71",
          5040 => x"2a",
          5041 => x"53",
          5042 => x"34",
          5043 => x"34",
          5044 => x"08",
          5045 => x"33",
          5046 => x"71",
          5047 => x"83",
          5048 => x"59",
          5049 => x"05",
          5050 => x"83",
          5051 => x"88",
          5052 => x"88",
          5053 => x"56",
          5054 => x"13",
          5055 => x"13",
          5056 => x"90",
          5057 => x"11",
          5058 => x"33",
          5059 => x"07",
          5060 => x"0c",
          5061 => x"3d",
          5062 => x"3d",
          5063 => x"b6",
          5064 => x"83",
          5065 => x"ff",
          5066 => x"53",
          5067 => x"a7",
          5068 => x"90",
          5069 => x"2b",
          5070 => x"11",
          5071 => x"33",
          5072 => x"71",
          5073 => x"75",
          5074 => x"81",
          5075 => x"98",
          5076 => x"2b",
          5077 => x"40",
          5078 => x"58",
          5079 => x"72",
          5080 => x"38",
          5081 => x"52",
          5082 => x"9d",
          5083 => x"39",
          5084 => x"85",
          5085 => x"8b",
          5086 => x"2b",
          5087 => x"79",
          5088 => x"51",
          5089 => x"76",
          5090 => x"75",
          5091 => x"56",
          5092 => x"34",
          5093 => x"08",
          5094 => x"12",
          5095 => x"33",
          5096 => x"07",
          5097 => x"54",
          5098 => x"53",
          5099 => x"34",
          5100 => x"34",
          5101 => x"08",
          5102 => x"0b",
          5103 => x"80",
          5104 => x"34",
          5105 => x"08",
          5106 => x"14",
          5107 => x"14",
          5108 => x"90",
          5109 => x"33",
          5110 => x"71",
          5111 => x"70",
          5112 => x"07",
          5113 => x"53",
          5114 => x"54",
          5115 => x"72",
          5116 => x"8b",
          5117 => x"ff",
          5118 => x"52",
          5119 => x"08",
          5120 => x"f2",
          5121 => x"2e",
          5122 => x"51",
          5123 => x"83",
          5124 => x"f5",
          5125 => x"7e",
          5126 => x"e2",
          5127 => x"98",
          5128 => x"ff",
          5129 => x"90",
          5130 => x"33",
          5131 => x"71",
          5132 => x"70",
          5133 => x"58",
          5134 => x"ff",
          5135 => x"2e",
          5136 => x"75",
          5137 => x"70",
          5138 => x"33",
          5139 => x"07",
          5140 => x"ff",
          5141 => x"70",
          5142 => x"06",
          5143 => x"52",
          5144 => x"59",
          5145 => x"27",
          5146 => x"80",
          5147 => x"75",
          5148 => x"84",
          5149 => x"16",
          5150 => x"2b",
          5151 => x"75",
          5152 => x"81",
          5153 => x"85",
          5154 => x"59",
          5155 => x"83",
          5156 => x"90",
          5157 => x"33",
          5158 => x"71",
          5159 => x"70",
          5160 => x"06",
          5161 => x"56",
          5162 => x"75",
          5163 => x"81",
          5164 => x"79",
          5165 => x"cc",
          5166 => x"74",
          5167 => x"c4",
          5168 => x"2e",
          5169 => x"89",
          5170 => x"f8",
          5171 => x"ac",
          5172 => x"80",
          5173 => x"75",
          5174 => x"3f",
          5175 => x"08",
          5176 => x"11",
          5177 => x"33",
          5178 => x"71",
          5179 => x"53",
          5180 => x"74",
          5181 => x"70",
          5182 => x"06",
          5183 => x"5c",
          5184 => x"78",
          5185 => x"76",
          5186 => x"57",
          5187 => x"34",
          5188 => x"08",
          5189 => x"71",
          5190 => x"86",
          5191 => x"12",
          5192 => x"2b",
          5193 => x"2a",
          5194 => x"53",
          5195 => x"73",
          5196 => x"75",
          5197 => x"82",
          5198 => x"70",
          5199 => x"33",
          5200 => x"71",
          5201 => x"83",
          5202 => x"5d",
          5203 => x"05",
          5204 => x"15",
          5205 => x"15",
          5206 => x"90",
          5207 => x"71",
          5208 => x"33",
          5209 => x"71",
          5210 => x"70",
          5211 => x"5a",
          5212 => x"54",
          5213 => x"34",
          5214 => x"34",
          5215 => x"08",
          5216 => x"54",
          5217 => x"98",
          5218 => x"0d",
          5219 => x"0d",
          5220 => x"b6",
          5221 => x"38",
          5222 => x"71",
          5223 => x"2e",
          5224 => x"51",
          5225 => x"82",
          5226 => x"53",
          5227 => x"98",
          5228 => x"0d",
          5229 => x"0d",
          5230 => x"5c",
          5231 => x"40",
          5232 => x"08",
          5233 => x"81",
          5234 => x"f4",
          5235 => x"8e",
          5236 => x"ff",
          5237 => x"b6",
          5238 => x"83",
          5239 => x"8b",
          5240 => x"fc",
          5241 => x"54",
          5242 => x"7e",
          5243 => x"3f",
          5244 => x"08",
          5245 => x"06",
          5246 => x"08",
          5247 => x"83",
          5248 => x"ff",
          5249 => x"83",
          5250 => x"70",
          5251 => x"33",
          5252 => x"07",
          5253 => x"70",
          5254 => x"06",
          5255 => x"fc",
          5256 => x"29",
          5257 => x"81",
          5258 => x"88",
          5259 => x"90",
          5260 => x"4e",
          5261 => x"52",
          5262 => x"41",
          5263 => x"5b",
          5264 => x"8f",
          5265 => x"ff",
          5266 => x"31",
          5267 => x"ff",
          5268 => x"82",
          5269 => x"17",
          5270 => x"2b",
          5271 => x"29",
          5272 => x"81",
          5273 => x"98",
          5274 => x"2b",
          5275 => x"45",
          5276 => x"73",
          5277 => x"38",
          5278 => x"70",
          5279 => x"06",
          5280 => x"7b",
          5281 => x"38",
          5282 => x"73",
          5283 => x"81",
          5284 => x"78",
          5285 => x"3f",
          5286 => x"ff",
          5287 => x"e5",
          5288 => x"38",
          5289 => x"89",
          5290 => x"f6",
          5291 => x"a5",
          5292 => x"55",
          5293 => x"80",
          5294 => x"1d",
          5295 => x"83",
          5296 => x"88",
          5297 => x"57",
          5298 => x"3f",
          5299 => x"51",
          5300 => x"82",
          5301 => x"83",
          5302 => x"7e",
          5303 => x"70",
          5304 => x"b6",
          5305 => x"84",
          5306 => x"59",
          5307 => x"3f",
          5308 => x"08",
          5309 => x"75",
          5310 => x"06",
          5311 => x"85",
          5312 => x"54",
          5313 => x"80",
          5314 => x"51",
          5315 => x"82",
          5316 => x"1d",
          5317 => x"83",
          5318 => x"88",
          5319 => x"43",
          5320 => x"3f",
          5321 => x"51",
          5322 => x"82",
          5323 => x"83",
          5324 => x"7e",
          5325 => x"70",
          5326 => x"b6",
          5327 => x"84",
          5328 => x"59",
          5329 => x"3f",
          5330 => x"08",
          5331 => x"60",
          5332 => x"55",
          5333 => x"ff",
          5334 => x"a9",
          5335 => x"52",
          5336 => x"3f",
          5337 => x"08",
          5338 => x"98",
          5339 => x"93",
          5340 => x"73",
          5341 => x"98",
          5342 => x"96",
          5343 => x"51",
          5344 => x"7a",
          5345 => x"27",
          5346 => x"53",
          5347 => x"51",
          5348 => x"7a",
          5349 => x"82",
          5350 => x"05",
          5351 => x"f6",
          5352 => x"54",
          5353 => x"98",
          5354 => x"0d",
          5355 => x"0d",
          5356 => x"70",
          5357 => x"d5",
          5358 => x"98",
          5359 => x"b6",
          5360 => x"2e",
          5361 => x"53",
          5362 => x"b6",
          5363 => x"ff",
          5364 => x"74",
          5365 => x"0c",
          5366 => x"04",
          5367 => x"02",
          5368 => x"51",
          5369 => x"72",
          5370 => x"82",
          5371 => x"33",
          5372 => x"b6",
          5373 => x"3d",
          5374 => x"3d",
          5375 => x"05",
          5376 => x"05",
          5377 => x"56",
          5378 => x"72",
          5379 => x"e0",
          5380 => x"2b",
          5381 => x"8c",
          5382 => x"88",
          5383 => x"2e",
          5384 => x"88",
          5385 => x"0c",
          5386 => x"8c",
          5387 => x"71",
          5388 => x"87",
          5389 => x"0c",
          5390 => x"08",
          5391 => x"51",
          5392 => x"2e",
          5393 => x"c0",
          5394 => x"51",
          5395 => x"71",
          5396 => x"80",
          5397 => x"92",
          5398 => x"98",
          5399 => x"70",
          5400 => x"38",
          5401 => x"94",
          5402 => x"b6",
          5403 => x"51",
          5404 => x"98",
          5405 => x"0d",
          5406 => x"0d",
          5407 => x"02",
          5408 => x"05",
          5409 => x"58",
          5410 => x"52",
          5411 => x"3f",
          5412 => x"08",
          5413 => x"54",
          5414 => x"be",
          5415 => x"75",
          5416 => x"c0",
          5417 => x"87",
          5418 => x"12",
          5419 => x"84",
          5420 => x"40",
          5421 => x"85",
          5422 => x"98",
          5423 => x"7d",
          5424 => x"0c",
          5425 => x"85",
          5426 => x"06",
          5427 => x"71",
          5428 => x"38",
          5429 => x"71",
          5430 => x"05",
          5431 => x"19",
          5432 => x"a2",
          5433 => x"71",
          5434 => x"38",
          5435 => x"83",
          5436 => x"38",
          5437 => x"8a",
          5438 => x"98",
          5439 => x"71",
          5440 => x"c0",
          5441 => x"52",
          5442 => x"87",
          5443 => x"80",
          5444 => x"81",
          5445 => x"c0",
          5446 => x"53",
          5447 => x"82",
          5448 => x"71",
          5449 => x"1a",
          5450 => x"84",
          5451 => x"19",
          5452 => x"06",
          5453 => x"79",
          5454 => x"38",
          5455 => x"80",
          5456 => x"87",
          5457 => x"26",
          5458 => x"73",
          5459 => x"06",
          5460 => x"2e",
          5461 => x"52",
          5462 => x"82",
          5463 => x"8f",
          5464 => x"f3",
          5465 => x"62",
          5466 => x"05",
          5467 => x"57",
          5468 => x"83",
          5469 => x"52",
          5470 => x"3f",
          5471 => x"08",
          5472 => x"54",
          5473 => x"2e",
          5474 => x"81",
          5475 => x"74",
          5476 => x"c0",
          5477 => x"87",
          5478 => x"12",
          5479 => x"84",
          5480 => x"5f",
          5481 => x"0b",
          5482 => x"8c",
          5483 => x"0c",
          5484 => x"80",
          5485 => x"70",
          5486 => x"81",
          5487 => x"54",
          5488 => x"8c",
          5489 => x"81",
          5490 => x"7c",
          5491 => x"58",
          5492 => x"70",
          5493 => x"52",
          5494 => x"8a",
          5495 => x"98",
          5496 => x"71",
          5497 => x"c0",
          5498 => x"52",
          5499 => x"87",
          5500 => x"80",
          5501 => x"81",
          5502 => x"c0",
          5503 => x"53",
          5504 => x"82",
          5505 => x"71",
          5506 => x"19",
          5507 => x"81",
          5508 => x"ff",
          5509 => x"19",
          5510 => x"78",
          5511 => x"38",
          5512 => x"80",
          5513 => x"87",
          5514 => x"26",
          5515 => x"73",
          5516 => x"06",
          5517 => x"2e",
          5518 => x"52",
          5519 => x"82",
          5520 => x"8f",
          5521 => x"fa",
          5522 => x"02",
          5523 => x"05",
          5524 => x"05",
          5525 => x"71",
          5526 => x"57",
          5527 => x"82",
          5528 => x"81",
          5529 => x"54",
          5530 => x"38",
          5531 => x"c0",
          5532 => x"81",
          5533 => x"2e",
          5534 => x"71",
          5535 => x"38",
          5536 => x"87",
          5537 => x"11",
          5538 => x"80",
          5539 => x"80",
          5540 => x"83",
          5541 => x"38",
          5542 => x"72",
          5543 => x"2a",
          5544 => x"51",
          5545 => x"80",
          5546 => x"87",
          5547 => x"08",
          5548 => x"38",
          5549 => x"8c",
          5550 => x"96",
          5551 => x"0c",
          5552 => x"8c",
          5553 => x"08",
          5554 => x"51",
          5555 => x"38",
          5556 => x"56",
          5557 => x"80",
          5558 => x"85",
          5559 => x"77",
          5560 => x"83",
          5561 => x"75",
          5562 => x"b6",
          5563 => x"3d",
          5564 => x"3d",
          5565 => x"11",
          5566 => x"71",
          5567 => x"82",
          5568 => x"53",
          5569 => x"0d",
          5570 => x"0d",
          5571 => x"33",
          5572 => x"71",
          5573 => x"88",
          5574 => x"14",
          5575 => x"07",
          5576 => x"33",
          5577 => x"b6",
          5578 => x"53",
          5579 => x"52",
          5580 => x"04",
          5581 => x"73",
          5582 => x"92",
          5583 => x"52",
          5584 => x"81",
          5585 => x"70",
          5586 => x"70",
          5587 => x"3d",
          5588 => x"3d",
          5589 => x"52",
          5590 => x"70",
          5591 => x"34",
          5592 => x"51",
          5593 => x"81",
          5594 => x"70",
          5595 => x"70",
          5596 => x"05",
          5597 => x"88",
          5598 => x"72",
          5599 => x"0d",
          5600 => x"0d",
          5601 => x"54",
          5602 => x"80",
          5603 => x"71",
          5604 => x"53",
          5605 => x"81",
          5606 => x"ff",
          5607 => x"39",
          5608 => x"04",
          5609 => x"75",
          5610 => x"52",
          5611 => x"70",
          5612 => x"34",
          5613 => x"70",
          5614 => x"3d",
          5615 => x"3d",
          5616 => x"79",
          5617 => x"74",
          5618 => x"56",
          5619 => x"81",
          5620 => x"71",
          5621 => x"16",
          5622 => x"52",
          5623 => x"86",
          5624 => x"2e",
          5625 => x"82",
          5626 => x"86",
          5627 => x"fe",
          5628 => x"76",
          5629 => x"39",
          5630 => x"8a",
          5631 => x"51",
          5632 => x"71",
          5633 => x"33",
          5634 => x"0c",
          5635 => x"04",
          5636 => x"b6",
          5637 => x"80",
          5638 => x"98",
          5639 => x"3d",
          5640 => x"80",
          5641 => x"33",
          5642 => x"7a",
          5643 => x"38",
          5644 => x"16",
          5645 => x"16",
          5646 => x"17",
          5647 => x"fa",
          5648 => x"b6",
          5649 => x"2e",
          5650 => x"b7",
          5651 => x"98",
          5652 => x"34",
          5653 => x"70",
          5654 => x"31",
          5655 => x"59",
          5656 => x"77",
          5657 => x"82",
          5658 => x"74",
          5659 => x"81",
          5660 => x"81",
          5661 => x"53",
          5662 => x"16",
          5663 => x"e3",
          5664 => x"81",
          5665 => x"b6",
          5666 => x"3d",
          5667 => x"3d",
          5668 => x"56",
          5669 => x"74",
          5670 => x"2e",
          5671 => x"51",
          5672 => x"82",
          5673 => x"57",
          5674 => x"08",
          5675 => x"54",
          5676 => x"16",
          5677 => x"33",
          5678 => x"3f",
          5679 => x"08",
          5680 => x"38",
          5681 => x"57",
          5682 => x"0c",
          5683 => x"98",
          5684 => x"0d",
          5685 => x"0d",
          5686 => x"57",
          5687 => x"82",
          5688 => x"58",
          5689 => x"08",
          5690 => x"76",
          5691 => x"83",
          5692 => x"06",
          5693 => x"84",
          5694 => x"78",
          5695 => x"81",
          5696 => x"38",
          5697 => x"82",
          5698 => x"52",
          5699 => x"52",
          5700 => x"3f",
          5701 => x"52",
          5702 => x"51",
          5703 => x"84",
          5704 => x"d2",
          5705 => x"fc",
          5706 => x"8a",
          5707 => x"52",
          5708 => x"51",
          5709 => x"90",
          5710 => x"84",
          5711 => x"fc",
          5712 => x"17",
          5713 => x"a0",
          5714 => x"86",
          5715 => x"08",
          5716 => x"b0",
          5717 => x"55",
          5718 => x"81",
          5719 => x"f8",
          5720 => x"84",
          5721 => x"53",
          5722 => x"17",
          5723 => x"d7",
          5724 => x"98",
          5725 => x"83",
          5726 => x"77",
          5727 => x"0c",
          5728 => x"04",
          5729 => x"77",
          5730 => x"12",
          5731 => x"55",
          5732 => x"56",
          5733 => x"8d",
          5734 => x"22",
          5735 => x"ac",
          5736 => x"57",
          5737 => x"b6",
          5738 => x"3d",
          5739 => x"3d",
          5740 => x"70",
          5741 => x"57",
          5742 => x"81",
          5743 => x"98",
          5744 => x"81",
          5745 => x"74",
          5746 => x"72",
          5747 => x"f5",
          5748 => x"24",
          5749 => x"81",
          5750 => x"81",
          5751 => x"83",
          5752 => x"38",
          5753 => x"76",
          5754 => x"70",
          5755 => x"16",
          5756 => x"74",
          5757 => x"96",
          5758 => x"98",
          5759 => x"38",
          5760 => x"06",
          5761 => x"33",
          5762 => x"89",
          5763 => x"08",
          5764 => x"54",
          5765 => x"fc",
          5766 => x"b6",
          5767 => x"fe",
          5768 => x"ff",
          5769 => x"11",
          5770 => x"2b",
          5771 => x"81",
          5772 => x"2a",
          5773 => x"51",
          5774 => x"e2",
          5775 => x"ff",
          5776 => x"da",
          5777 => x"2a",
          5778 => x"05",
          5779 => x"fc",
          5780 => x"b6",
          5781 => x"c6",
          5782 => x"83",
          5783 => x"05",
          5784 => x"f9",
          5785 => x"b6",
          5786 => x"ff",
          5787 => x"ae",
          5788 => x"2a",
          5789 => x"05",
          5790 => x"fc",
          5791 => x"b6",
          5792 => x"38",
          5793 => x"83",
          5794 => x"05",
          5795 => x"f8",
          5796 => x"b6",
          5797 => x"0a",
          5798 => x"39",
          5799 => x"82",
          5800 => x"89",
          5801 => x"f8",
          5802 => x"7c",
          5803 => x"56",
          5804 => x"77",
          5805 => x"38",
          5806 => x"08",
          5807 => x"38",
          5808 => x"72",
          5809 => x"9d",
          5810 => x"24",
          5811 => x"81",
          5812 => x"82",
          5813 => x"83",
          5814 => x"38",
          5815 => x"76",
          5816 => x"70",
          5817 => x"18",
          5818 => x"76",
          5819 => x"9e",
          5820 => x"98",
          5821 => x"b6",
          5822 => x"d9",
          5823 => x"ff",
          5824 => x"05",
          5825 => x"81",
          5826 => x"54",
          5827 => x"80",
          5828 => x"77",
          5829 => x"f0",
          5830 => x"8f",
          5831 => x"51",
          5832 => x"34",
          5833 => x"17",
          5834 => x"2a",
          5835 => x"05",
          5836 => x"fa",
          5837 => x"b6",
          5838 => x"82",
          5839 => x"81",
          5840 => x"83",
          5841 => x"b4",
          5842 => x"2a",
          5843 => x"8f",
          5844 => x"2a",
          5845 => x"f0",
          5846 => x"06",
          5847 => x"72",
          5848 => x"ec",
          5849 => x"2a",
          5850 => x"05",
          5851 => x"fa",
          5852 => x"b6",
          5853 => x"82",
          5854 => x"80",
          5855 => x"83",
          5856 => x"52",
          5857 => x"fe",
          5858 => x"b4",
          5859 => x"a4",
          5860 => x"76",
          5861 => x"17",
          5862 => x"75",
          5863 => x"3f",
          5864 => x"08",
          5865 => x"98",
          5866 => x"77",
          5867 => x"77",
          5868 => x"fc",
          5869 => x"b4",
          5870 => x"51",
          5871 => x"c9",
          5872 => x"98",
          5873 => x"06",
          5874 => x"72",
          5875 => x"3f",
          5876 => x"17",
          5877 => x"b6",
          5878 => x"3d",
          5879 => x"3d",
          5880 => x"7e",
          5881 => x"56",
          5882 => x"75",
          5883 => x"74",
          5884 => x"27",
          5885 => x"80",
          5886 => x"ff",
          5887 => x"75",
          5888 => x"3f",
          5889 => x"08",
          5890 => x"98",
          5891 => x"38",
          5892 => x"54",
          5893 => x"81",
          5894 => x"39",
          5895 => x"08",
          5896 => x"39",
          5897 => x"51",
          5898 => x"82",
          5899 => x"58",
          5900 => x"08",
          5901 => x"c7",
          5902 => x"98",
          5903 => x"d2",
          5904 => x"98",
          5905 => x"cf",
          5906 => x"74",
          5907 => x"fc",
          5908 => x"b6",
          5909 => x"38",
          5910 => x"fe",
          5911 => x"08",
          5912 => x"74",
          5913 => x"38",
          5914 => x"17",
          5915 => x"33",
          5916 => x"73",
          5917 => x"77",
          5918 => x"26",
          5919 => x"80",
          5920 => x"b6",
          5921 => x"3d",
          5922 => x"3d",
          5923 => x"71",
          5924 => x"5b",
          5925 => x"8c",
          5926 => x"77",
          5927 => x"38",
          5928 => x"78",
          5929 => x"81",
          5930 => x"79",
          5931 => x"f9",
          5932 => x"55",
          5933 => x"98",
          5934 => x"e0",
          5935 => x"98",
          5936 => x"b6",
          5937 => x"2e",
          5938 => x"98",
          5939 => x"b6",
          5940 => x"82",
          5941 => x"58",
          5942 => x"70",
          5943 => x"80",
          5944 => x"38",
          5945 => x"09",
          5946 => x"e2",
          5947 => x"56",
          5948 => x"76",
          5949 => x"82",
          5950 => x"7a",
          5951 => x"3f",
          5952 => x"b6",
          5953 => x"2e",
          5954 => x"86",
          5955 => x"98",
          5956 => x"b6",
          5957 => x"70",
          5958 => x"07",
          5959 => x"7c",
          5960 => x"98",
          5961 => x"51",
          5962 => x"81",
          5963 => x"b6",
          5964 => x"2e",
          5965 => x"17",
          5966 => x"74",
          5967 => x"73",
          5968 => x"27",
          5969 => x"58",
          5970 => x"80",
          5971 => x"56",
          5972 => x"98",
          5973 => x"26",
          5974 => x"56",
          5975 => x"81",
          5976 => x"52",
          5977 => x"c6",
          5978 => x"98",
          5979 => x"b8",
          5980 => x"82",
          5981 => x"81",
          5982 => x"06",
          5983 => x"b6",
          5984 => x"82",
          5985 => x"09",
          5986 => x"72",
          5987 => x"70",
          5988 => x"51",
          5989 => x"80",
          5990 => x"78",
          5991 => x"06",
          5992 => x"73",
          5993 => x"39",
          5994 => x"52",
          5995 => x"f7",
          5996 => x"98",
          5997 => x"98",
          5998 => x"82",
          5999 => x"07",
          6000 => x"55",
          6001 => x"2e",
          6002 => x"80",
          6003 => x"75",
          6004 => x"76",
          6005 => x"3f",
          6006 => x"08",
          6007 => x"38",
          6008 => x"0c",
          6009 => x"fe",
          6010 => x"08",
          6011 => x"74",
          6012 => x"ff",
          6013 => x"0c",
          6014 => x"81",
          6015 => x"84",
          6016 => x"39",
          6017 => x"81",
          6018 => x"8c",
          6019 => x"8c",
          6020 => x"98",
          6021 => x"39",
          6022 => x"55",
          6023 => x"98",
          6024 => x"0d",
          6025 => x"0d",
          6026 => x"55",
          6027 => x"82",
          6028 => x"58",
          6029 => x"b6",
          6030 => x"d8",
          6031 => x"74",
          6032 => x"3f",
          6033 => x"08",
          6034 => x"08",
          6035 => x"59",
          6036 => x"77",
          6037 => x"70",
          6038 => x"c8",
          6039 => x"84",
          6040 => x"56",
          6041 => x"58",
          6042 => x"97",
          6043 => x"75",
          6044 => x"52",
          6045 => x"51",
          6046 => x"82",
          6047 => x"80",
          6048 => x"8a",
          6049 => x"32",
          6050 => x"72",
          6051 => x"2a",
          6052 => x"56",
          6053 => x"98",
          6054 => x"0d",
          6055 => x"0d",
          6056 => x"08",
          6057 => x"74",
          6058 => x"26",
          6059 => x"74",
          6060 => x"72",
          6061 => x"74",
          6062 => x"88",
          6063 => x"73",
          6064 => x"33",
          6065 => x"27",
          6066 => x"16",
          6067 => x"9b",
          6068 => x"2a",
          6069 => x"88",
          6070 => x"58",
          6071 => x"80",
          6072 => x"16",
          6073 => x"0c",
          6074 => x"8a",
          6075 => x"89",
          6076 => x"72",
          6077 => x"38",
          6078 => x"51",
          6079 => x"82",
          6080 => x"54",
          6081 => x"08",
          6082 => x"38",
          6083 => x"b6",
          6084 => x"8b",
          6085 => x"08",
          6086 => x"08",
          6087 => x"82",
          6088 => x"74",
          6089 => x"cb",
          6090 => x"75",
          6091 => x"3f",
          6092 => x"08",
          6093 => x"73",
          6094 => x"98",
          6095 => x"82",
          6096 => x"2e",
          6097 => x"39",
          6098 => x"39",
          6099 => x"13",
          6100 => x"74",
          6101 => x"16",
          6102 => x"18",
          6103 => x"77",
          6104 => x"0c",
          6105 => x"04",
          6106 => x"7a",
          6107 => x"12",
          6108 => x"59",
          6109 => x"80",
          6110 => x"86",
          6111 => x"98",
          6112 => x"14",
          6113 => x"55",
          6114 => x"81",
          6115 => x"83",
          6116 => x"77",
          6117 => x"81",
          6118 => x"0c",
          6119 => x"55",
          6120 => x"76",
          6121 => x"17",
          6122 => x"74",
          6123 => x"9b",
          6124 => x"39",
          6125 => x"ff",
          6126 => x"2a",
          6127 => x"81",
          6128 => x"52",
          6129 => x"e6",
          6130 => x"98",
          6131 => x"55",
          6132 => x"b6",
          6133 => x"80",
          6134 => x"55",
          6135 => x"08",
          6136 => x"f4",
          6137 => x"08",
          6138 => x"08",
          6139 => x"38",
          6140 => x"77",
          6141 => x"84",
          6142 => x"39",
          6143 => x"52",
          6144 => x"86",
          6145 => x"98",
          6146 => x"55",
          6147 => x"08",
          6148 => x"c4",
          6149 => x"82",
          6150 => x"81",
          6151 => x"81",
          6152 => x"98",
          6153 => x"b0",
          6154 => x"98",
          6155 => x"51",
          6156 => x"82",
          6157 => x"a0",
          6158 => x"15",
          6159 => x"75",
          6160 => x"3f",
          6161 => x"08",
          6162 => x"76",
          6163 => x"77",
          6164 => x"9c",
          6165 => x"55",
          6166 => x"98",
          6167 => x"0d",
          6168 => x"0d",
          6169 => x"08",
          6170 => x"80",
          6171 => x"fc",
          6172 => x"b6",
          6173 => x"82",
          6174 => x"80",
          6175 => x"b6",
          6176 => x"98",
          6177 => x"78",
          6178 => x"3f",
          6179 => x"08",
          6180 => x"98",
          6181 => x"38",
          6182 => x"08",
          6183 => x"70",
          6184 => x"58",
          6185 => x"2e",
          6186 => x"83",
          6187 => x"82",
          6188 => x"55",
          6189 => x"81",
          6190 => x"07",
          6191 => x"2e",
          6192 => x"16",
          6193 => x"2e",
          6194 => x"88",
          6195 => x"82",
          6196 => x"56",
          6197 => x"51",
          6198 => x"82",
          6199 => x"54",
          6200 => x"08",
          6201 => x"9b",
          6202 => x"2e",
          6203 => x"83",
          6204 => x"73",
          6205 => x"0c",
          6206 => x"04",
          6207 => x"76",
          6208 => x"54",
          6209 => x"82",
          6210 => x"83",
          6211 => x"76",
          6212 => x"53",
          6213 => x"2e",
          6214 => x"90",
          6215 => x"51",
          6216 => x"82",
          6217 => x"90",
          6218 => x"53",
          6219 => x"98",
          6220 => x"0d",
          6221 => x"0d",
          6222 => x"83",
          6223 => x"54",
          6224 => x"55",
          6225 => x"3f",
          6226 => x"51",
          6227 => x"2e",
          6228 => x"8b",
          6229 => x"2a",
          6230 => x"51",
          6231 => x"86",
          6232 => x"f7",
          6233 => x"7d",
          6234 => x"75",
          6235 => x"98",
          6236 => x"2e",
          6237 => x"98",
          6238 => x"78",
          6239 => x"3f",
          6240 => x"08",
          6241 => x"98",
          6242 => x"38",
          6243 => x"70",
          6244 => x"73",
          6245 => x"58",
          6246 => x"8b",
          6247 => x"bf",
          6248 => x"ff",
          6249 => x"53",
          6250 => x"34",
          6251 => x"08",
          6252 => x"e5",
          6253 => x"81",
          6254 => x"2e",
          6255 => x"70",
          6256 => x"57",
          6257 => x"9e",
          6258 => x"2e",
          6259 => x"b6",
          6260 => x"df",
          6261 => x"72",
          6262 => x"81",
          6263 => x"76",
          6264 => x"2e",
          6265 => x"52",
          6266 => x"fc",
          6267 => x"98",
          6268 => x"b6",
          6269 => x"38",
          6270 => x"fe",
          6271 => x"39",
          6272 => x"16",
          6273 => x"b6",
          6274 => x"3d",
          6275 => x"3d",
          6276 => x"08",
          6277 => x"52",
          6278 => x"c5",
          6279 => x"98",
          6280 => x"b6",
          6281 => x"38",
          6282 => x"52",
          6283 => x"de",
          6284 => x"98",
          6285 => x"b6",
          6286 => x"38",
          6287 => x"b6",
          6288 => x"9c",
          6289 => x"ea",
          6290 => x"53",
          6291 => x"9c",
          6292 => x"ea",
          6293 => x"0b",
          6294 => x"74",
          6295 => x"0c",
          6296 => x"04",
          6297 => x"75",
          6298 => x"12",
          6299 => x"53",
          6300 => x"9a",
          6301 => x"98",
          6302 => x"9c",
          6303 => x"e5",
          6304 => x"0b",
          6305 => x"85",
          6306 => x"fa",
          6307 => x"7a",
          6308 => x"0b",
          6309 => x"98",
          6310 => x"2e",
          6311 => x"80",
          6312 => x"55",
          6313 => x"17",
          6314 => x"33",
          6315 => x"51",
          6316 => x"2e",
          6317 => x"85",
          6318 => x"06",
          6319 => x"e5",
          6320 => x"2e",
          6321 => x"8b",
          6322 => x"70",
          6323 => x"34",
          6324 => x"71",
          6325 => x"05",
          6326 => x"15",
          6327 => x"27",
          6328 => x"15",
          6329 => x"80",
          6330 => x"34",
          6331 => x"52",
          6332 => x"88",
          6333 => x"17",
          6334 => x"52",
          6335 => x"3f",
          6336 => x"08",
          6337 => x"12",
          6338 => x"3f",
          6339 => x"08",
          6340 => x"98",
          6341 => x"da",
          6342 => x"98",
          6343 => x"23",
          6344 => x"04",
          6345 => x"7f",
          6346 => x"5b",
          6347 => x"33",
          6348 => x"73",
          6349 => x"38",
          6350 => x"80",
          6351 => x"38",
          6352 => x"8c",
          6353 => x"08",
          6354 => x"aa",
          6355 => x"41",
          6356 => x"33",
          6357 => x"73",
          6358 => x"81",
          6359 => x"81",
          6360 => x"dc",
          6361 => x"70",
          6362 => x"07",
          6363 => x"73",
          6364 => x"88",
          6365 => x"70",
          6366 => x"73",
          6367 => x"38",
          6368 => x"ab",
          6369 => x"52",
          6370 => x"91",
          6371 => x"98",
          6372 => x"98",
          6373 => x"61",
          6374 => x"5a",
          6375 => x"a0",
          6376 => x"e7",
          6377 => x"70",
          6378 => x"79",
          6379 => x"73",
          6380 => x"81",
          6381 => x"38",
          6382 => x"33",
          6383 => x"ae",
          6384 => x"70",
          6385 => x"82",
          6386 => x"51",
          6387 => x"54",
          6388 => x"79",
          6389 => x"74",
          6390 => x"57",
          6391 => x"af",
          6392 => x"70",
          6393 => x"51",
          6394 => x"dc",
          6395 => x"73",
          6396 => x"38",
          6397 => x"82",
          6398 => x"19",
          6399 => x"54",
          6400 => x"82",
          6401 => x"54",
          6402 => x"78",
          6403 => x"81",
          6404 => x"54",
          6405 => x"81",
          6406 => x"af",
          6407 => x"77",
          6408 => x"70",
          6409 => x"25",
          6410 => x"07",
          6411 => x"51",
          6412 => x"2e",
          6413 => x"39",
          6414 => x"80",
          6415 => x"33",
          6416 => x"73",
          6417 => x"81",
          6418 => x"81",
          6419 => x"dc",
          6420 => x"70",
          6421 => x"07",
          6422 => x"73",
          6423 => x"b5",
          6424 => x"2e",
          6425 => x"83",
          6426 => x"76",
          6427 => x"07",
          6428 => x"2e",
          6429 => x"8b",
          6430 => x"77",
          6431 => x"30",
          6432 => x"71",
          6433 => x"53",
          6434 => x"55",
          6435 => x"38",
          6436 => x"5c",
          6437 => x"75",
          6438 => x"73",
          6439 => x"38",
          6440 => x"06",
          6441 => x"11",
          6442 => x"75",
          6443 => x"3f",
          6444 => x"08",
          6445 => x"38",
          6446 => x"33",
          6447 => x"54",
          6448 => x"e6",
          6449 => x"b6",
          6450 => x"2e",
          6451 => x"ff",
          6452 => x"74",
          6453 => x"38",
          6454 => x"75",
          6455 => x"17",
          6456 => x"57",
          6457 => x"a7",
          6458 => x"82",
          6459 => x"e5",
          6460 => x"b6",
          6461 => x"38",
          6462 => x"54",
          6463 => x"89",
          6464 => x"70",
          6465 => x"57",
          6466 => x"54",
          6467 => x"81",
          6468 => x"f7",
          6469 => x"7e",
          6470 => x"2e",
          6471 => x"33",
          6472 => x"e5",
          6473 => x"06",
          6474 => x"7a",
          6475 => x"a0",
          6476 => x"38",
          6477 => x"55",
          6478 => x"84",
          6479 => x"39",
          6480 => x"8b",
          6481 => x"7b",
          6482 => x"7a",
          6483 => x"3f",
          6484 => x"08",
          6485 => x"98",
          6486 => x"38",
          6487 => x"52",
          6488 => x"aa",
          6489 => x"98",
          6490 => x"b6",
          6491 => x"c2",
          6492 => x"08",
          6493 => x"55",
          6494 => x"ff",
          6495 => x"15",
          6496 => x"54",
          6497 => x"34",
          6498 => x"70",
          6499 => x"81",
          6500 => x"58",
          6501 => x"8b",
          6502 => x"74",
          6503 => x"3f",
          6504 => x"08",
          6505 => x"38",
          6506 => x"51",
          6507 => x"ff",
          6508 => x"ab",
          6509 => x"55",
          6510 => x"bb",
          6511 => x"2e",
          6512 => x"80",
          6513 => x"85",
          6514 => x"06",
          6515 => x"58",
          6516 => x"80",
          6517 => x"75",
          6518 => x"73",
          6519 => x"b5",
          6520 => x"0b",
          6521 => x"80",
          6522 => x"39",
          6523 => x"54",
          6524 => x"85",
          6525 => x"75",
          6526 => x"81",
          6527 => x"73",
          6528 => x"1b",
          6529 => x"2a",
          6530 => x"51",
          6531 => x"80",
          6532 => x"90",
          6533 => x"ff",
          6534 => x"05",
          6535 => x"f5",
          6536 => x"b6",
          6537 => x"1c",
          6538 => x"39",
          6539 => x"98",
          6540 => x"0d",
          6541 => x"0d",
          6542 => x"7b",
          6543 => x"73",
          6544 => x"55",
          6545 => x"2e",
          6546 => x"75",
          6547 => x"57",
          6548 => x"26",
          6549 => x"ba",
          6550 => x"70",
          6551 => x"ba",
          6552 => x"06",
          6553 => x"73",
          6554 => x"70",
          6555 => x"51",
          6556 => x"89",
          6557 => x"82",
          6558 => x"ff",
          6559 => x"56",
          6560 => x"2e",
          6561 => x"80",
          6562 => x"d0",
          6563 => x"08",
          6564 => x"76",
          6565 => x"58",
          6566 => x"81",
          6567 => x"ff",
          6568 => x"53",
          6569 => x"26",
          6570 => x"13",
          6571 => x"06",
          6572 => x"9f",
          6573 => x"99",
          6574 => x"e0",
          6575 => x"ff",
          6576 => x"72",
          6577 => x"2a",
          6578 => x"72",
          6579 => x"06",
          6580 => x"ff",
          6581 => x"30",
          6582 => x"70",
          6583 => x"07",
          6584 => x"9f",
          6585 => x"54",
          6586 => x"80",
          6587 => x"81",
          6588 => x"59",
          6589 => x"25",
          6590 => x"8b",
          6591 => x"24",
          6592 => x"76",
          6593 => x"78",
          6594 => x"82",
          6595 => x"51",
          6596 => x"98",
          6597 => x"0d",
          6598 => x"0d",
          6599 => x"0b",
          6600 => x"ff",
          6601 => x"0c",
          6602 => x"51",
          6603 => x"84",
          6604 => x"98",
          6605 => x"38",
          6606 => x"51",
          6607 => x"82",
          6608 => x"83",
          6609 => x"54",
          6610 => x"82",
          6611 => x"09",
          6612 => x"e3",
          6613 => x"b4",
          6614 => x"57",
          6615 => x"2e",
          6616 => x"83",
          6617 => x"74",
          6618 => x"70",
          6619 => x"25",
          6620 => x"51",
          6621 => x"38",
          6622 => x"2e",
          6623 => x"b5",
          6624 => x"82",
          6625 => x"80",
          6626 => x"e0",
          6627 => x"b6",
          6628 => x"82",
          6629 => x"80",
          6630 => x"85",
          6631 => x"94",
          6632 => x"16",
          6633 => x"3f",
          6634 => x"08",
          6635 => x"98",
          6636 => x"83",
          6637 => x"74",
          6638 => x"0c",
          6639 => x"04",
          6640 => x"61",
          6641 => x"80",
          6642 => x"58",
          6643 => x"0c",
          6644 => x"e1",
          6645 => x"98",
          6646 => x"56",
          6647 => x"b6",
          6648 => x"86",
          6649 => x"b6",
          6650 => x"29",
          6651 => x"05",
          6652 => x"53",
          6653 => x"80",
          6654 => x"38",
          6655 => x"76",
          6656 => x"74",
          6657 => x"72",
          6658 => x"38",
          6659 => x"51",
          6660 => x"82",
          6661 => x"81",
          6662 => x"81",
          6663 => x"72",
          6664 => x"80",
          6665 => x"38",
          6666 => x"70",
          6667 => x"53",
          6668 => x"86",
          6669 => x"a7",
          6670 => x"34",
          6671 => x"34",
          6672 => x"14",
          6673 => x"b2",
          6674 => x"98",
          6675 => x"06",
          6676 => x"54",
          6677 => x"72",
          6678 => x"76",
          6679 => x"38",
          6680 => x"70",
          6681 => x"53",
          6682 => x"85",
          6683 => x"70",
          6684 => x"5b",
          6685 => x"82",
          6686 => x"81",
          6687 => x"76",
          6688 => x"81",
          6689 => x"38",
          6690 => x"56",
          6691 => x"83",
          6692 => x"70",
          6693 => x"80",
          6694 => x"83",
          6695 => x"dc",
          6696 => x"b6",
          6697 => x"76",
          6698 => x"05",
          6699 => x"16",
          6700 => x"56",
          6701 => x"d7",
          6702 => x"8d",
          6703 => x"72",
          6704 => x"54",
          6705 => x"57",
          6706 => x"95",
          6707 => x"73",
          6708 => x"3f",
          6709 => x"08",
          6710 => x"57",
          6711 => x"89",
          6712 => x"56",
          6713 => x"d7",
          6714 => x"76",
          6715 => x"f1",
          6716 => x"76",
          6717 => x"e9",
          6718 => x"51",
          6719 => x"82",
          6720 => x"83",
          6721 => x"53",
          6722 => x"2e",
          6723 => x"84",
          6724 => x"ca",
          6725 => x"da",
          6726 => x"98",
          6727 => x"ff",
          6728 => x"8d",
          6729 => x"14",
          6730 => x"3f",
          6731 => x"08",
          6732 => x"15",
          6733 => x"14",
          6734 => x"34",
          6735 => x"33",
          6736 => x"81",
          6737 => x"54",
          6738 => x"72",
          6739 => x"91",
          6740 => x"ff",
          6741 => x"29",
          6742 => x"33",
          6743 => x"72",
          6744 => x"72",
          6745 => x"38",
          6746 => x"06",
          6747 => x"2e",
          6748 => x"56",
          6749 => x"80",
          6750 => x"da",
          6751 => x"b6",
          6752 => x"82",
          6753 => x"88",
          6754 => x"8f",
          6755 => x"56",
          6756 => x"38",
          6757 => x"51",
          6758 => x"82",
          6759 => x"83",
          6760 => x"55",
          6761 => x"80",
          6762 => x"da",
          6763 => x"b6",
          6764 => x"80",
          6765 => x"da",
          6766 => x"b6",
          6767 => x"ff",
          6768 => x"8d",
          6769 => x"2e",
          6770 => x"88",
          6771 => x"14",
          6772 => x"05",
          6773 => x"75",
          6774 => x"38",
          6775 => x"52",
          6776 => x"51",
          6777 => x"3f",
          6778 => x"08",
          6779 => x"98",
          6780 => x"82",
          6781 => x"b6",
          6782 => x"ff",
          6783 => x"26",
          6784 => x"57",
          6785 => x"f5",
          6786 => x"82",
          6787 => x"f5",
          6788 => x"81",
          6789 => x"8d",
          6790 => x"2e",
          6791 => x"82",
          6792 => x"16",
          6793 => x"16",
          6794 => x"70",
          6795 => x"7a",
          6796 => x"0c",
          6797 => x"83",
          6798 => x"06",
          6799 => x"de",
          6800 => x"ae",
          6801 => x"98",
          6802 => x"ff",
          6803 => x"56",
          6804 => x"38",
          6805 => x"38",
          6806 => x"51",
          6807 => x"82",
          6808 => x"a8",
          6809 => x"82",
          6810 => x"39",
          6811 => x"80",
          6812 => x"38",
          6813 => x"15",
          6814 => x"53",
          6815 => x"8d",
          6816 => x"15",
          6817 => x"76",
          6818 => x"51",
          6819 => x"13",
          6820 => x"8d",
          6821 => x"15",
          6822 => x"c5",
          6823 => x"90",
          6824 => x"0b",
          6825 => x"ff",
          6826 => x"15",
          6827 => x"2e",
          6828 => x"81",
          6829 => x"e4",
          6830 => x"b6",
          6831 => x"98",
          6832 => x"ff",
          6833 => x"81",
          6834 => x"06",
          6835 => x"81",
          6836 => x"51",
          6837 => x"82",
          6838 => x"80",
          6839 => x"b6",
          6840 => x"15",
          6841 => x"14",
          6842 => x"3f",
          6843 => x"08",
          6844 => x"06",
          6845 => x"d4",
          6846 => x"81",
          6847 => x"38",
          6848 => x"d8",
          6849 => x"b6",
          6850 => x"8b",
          6851 => x"2e",
          6852 => x"b3",
          6853 => x"14",
          6854 => x"3f",
          6855 => x"08",
          6856 => x"e4",
          6857 => x"81",
          6858 => x"84",
          6859 => x"d7",
          6860 => x"b6",
          6861 => x"15",
          6862 => x"14",
          6863 => x"3f",
          6864 => x"08",
          6865 => x"76",
          6866 => x"cd",
          6867 => x"05",
          6868 => x"cd",
          6869 => x"86",
          6870 => x"0b",
          6871 => x"80",
          6872 => x"b6",
          6873 => x"3d",
          6874 => x"3d",
          6875 => x"89",
          6876 => x"2e",
          6877 => x"08",
          6878 => x"2e",
          6879 => x"33",
          6880 => x"2e",
          6881 => x"13",
          6882 => x"22",
          6883 => x"76",
          6884 => x"06",
          6885 => x"13",
          6886 => x"c0",
          6887 => x"98",
          6888 => x"52",
          6889 => x"71",
          6890 => x"55",
          6891 => x"53",
          6892 => x"0c",
          6893 => x"b6",
          6894 => x"3d",
          6895 => x"3d",
          6896 => x"05",
          6897 => x"89",
          6898 => x"52",
          6899 => x"3f",
          6900 => x"0b",
          6901 => x"08",
          6902 => x"82",
          6903 => x"84",
          6904 => x"d0",
          6905 => x"55",
          6906 => x"2e",
          6907 => x"74",
          6908 => x"73",
          6909 => x"38",
          6910 => x"78",
          6911 => x"54",
          6912 => x"92",
          6913 => x"89",
          6914 => x"84",
          6915 => x"b0",
          6916 => x"98",
          6917 => x"82",
          6918 => x"88",
          6919 => x"eb",
          6920 => x"02",
          6921 => x"e7",
          6922 => x"59",
          6923 => x"80",
          6924 => x"38",
          6925 => x"70",
          6926 => x"d0",
          6927 => x"3d",
          6928 => x"58",
          6929 => x"82",
          6930 => x"55",
          6931 => x"08",
          6932 => x"7a",
          6933 => x"8c",
          6934 => x"56",
          6935 => x"82",
          6936 => x"55",
          6937 => x"08",
          6938 => x"80",
          6939 => x"70",
          6940 => x"57",
          6941 => x"83",
          6942 => x"77",
          6943 => x"73",
          6944 => x"ab",
          6945 => x"2e",
          6946 => x"84",
          6947 => x"06",
          6948 => x"51",
          6949 => x"82",
          6950 => x"55",
          6951 => x"b2",
          6952 => x"06",
          6953 => x"b8",
          6954 => x"2a",
          6955 => x"51",
          6956 => x"2e",
          6957 => x"55",
          6958 => x"77",
          6959 => x"74",
          6960 => x"77",
          6961 => x"81",
          6962 => x"73",
          6963 => x"af",
          6964 => x"7a",
          6965 => x"3f",
          6966 => x"08",
          6967 => x"b2",
          6968 => x"8e",
          6969 => x"ea",
          6970 => x"a0",
          6971 => x"34",
          6972 => x"52",
          6973 => x"bd",
          6974 => x"62",
          6975 => x"d4",
          6976 => x"54",
          6977 => x"15",
          6978 => x"2e",
          6979 => x"7a",
          6980 => x"51",
          6981 => x"75",
          6982 => x"d4",
          6983 => x"be",
          6984 => x"98",
          6985 => x"b6",
          6986 => x"ca",
          6987 => x"74",
          6988 => x"02",
          6989 => x"70",
          6990 => x"81",
          6991 => x"56",
          6992 => x"86",
          6993 => x"82",
          6994 => x"81",
          6995 => x"06",
          6996 => x"80",
          6997 => x"75",
          6998 => x"73",
          6999 => x"38",
          7000 => x"92",
          7001 => x"7a",
          7002 => x"3f",
          7003 => x"08",
          7004 => x"8c",
          7005 => x"55",
          7006 => x"08",
          7007 => x"77",
          7008 => x"81",
          7009 => x"73",
          7010 => x"38",
          7011 => x"07",
          7012 => x"11",
          7013 => x"0c",
          7014 => x"0c",
          7015 => x"52",
          7016 => x"3f",
          7017 => x"08",
          7018 => x"08",
          7019 => x"63",
          7020 => x"5a",
          7021 => x"82",
          7022 => x"82",
          7023 => x"8c",
          7024 => x"7a",
          7025 => x"17",
          7026 => x"23",
          7027 => x"34",
          7028 => x"1a",
          7029 => x"9c",
          7030 => x"0b",
          7031 => x"77",
          7032 => x"81",
          7033 => x"73",
          7034 => x"8d",
          7035 => x"98",
          7036 => x"81",
          7037 => x"b6",
          7038 => x"1a",
          7039 => x"22",
          7040 => x"7b",
          7041 => x"a8",
          7042 => x"78",
          7043 => x"3f",
          7044 => x"08",
          7045 => x"98",
          7046 => x"83",
          7047 => x"82",
          7048 => x"ff",
          7049 => x"06",
          7050 => x"55",
          7051 => x"56",
          7052 => x"76",
          7053 => x"51",
          7054 => x"27",
          7055 => x"70",
          7056 => x"5a",
          7057 => x"76",
          7058 => x"74",
          7059 => x"83",
          7060 => x"73",
          7061 => x"38",
          7062 => x"51",
          7063 => x"82",
          7064 => x"85",
          7065 => x"8e",
          7066 => x"2a",
          7067 => x"08",
          7068 => x"0c",
          7069 => x"79",
          7070 => x"73",
          7071 => x"0c",
          7072 => x"04",
          7073 => x"60",
          7074 => x"40",
          7075 => x"80",
          7076 => x"3d",
          7077 => x"78",
          7078 => x"3f",
          7079 => x"08",
          7080 => x"98",
          7081 => x"91",
          7082 => x"74",
          7083 => x"38",
          7084 => x"c4",
          7085 => x"33",
          7086 => x"87",
          7087 => x"2e",
          7088 => x"95",
          7089 => x"91",
          7090 => x"56",
          7091 => x"81",
          7092 => x"34",
          7093 => x"a0",
          7094 => x"08",
          7095 => x"31",
          7096 => x"27",
          7097 => x"5c",
          7098 => x"82",
          7099 => x"19",
          7100 => x"ff",
          7101 => x"74",
          7102 => x"7e",
          7103 => x"ff",
          7104 => x"2a",
          7105 => x"79",
          7106 => x"87",
          7107 => x"08",
          7108 => x"98",
          7109 => x"78",
          7110 => x"3f",
          7111 => x"08",
          7112 => x"27",
          7113 => x"74",
          7114 => x"a3",
          7115 => x"1a",
          7116 => x"08",
          7117 => x"d4",
          7118 => x"b6",
          7119 => x"2e",
          7120 => x"82",
          7121 => x"1a",
          7122 => x"59",
          7123 => x"2e",
          7124 => x"77",
          7125 => x"11",
          7126 => x"55",
          7127 => x"85",
          7128 => x"31",
          7129 => x"76",
          7130 => x"81",
          7131 => x"ca",
          7132 => x"b6",
          7133 => x"d7",
          7134 => x"11",
          7135 => x"74",
          7136 => x"38",
          7137 => x"77",
          7138 => x"78",
          7139 => x"84",
          7140 => x"16",
          7141 => x"08",
          7142 => x"2b",
          7143 => x"cf",
          7144 => x"89",
          7145 => x"39",
          7146 => x"0c",
          7147 => x"83",
          7148 => x"80",
          7149 => x"55",
          7150 => x"83",
          7151 => x"9c",
          7152 => x"7e",
          7153 => x"3f",
          7154 => x"08",
          7155 => x"75",
          7156 => x"08",
          7157 => x"1f",
          7158 => x"7c",
          7159 => x"3f",
          7160 => x"7e",
          7161 => x"0c",
          7162 => x"1b",
          7163 => x"1c",
          7164 => x"fd",
          7165 => x"56",
          7166 => x"98",
          7167 => x"0d",
          7168 => x"0d",
          7169 => x"64",
          7170 => x"58",
          7171 => x"90",
          7172 => x"52",
          7173 => x"d2",
          7174 => x"98",
          7175 => x"b6",
          7176 => x"38",
          7177 => x"55",
          7178 => x"86",
          7179 => x"83",
          7180 => x"18",
          7181 => x"2a",
          7182 => x"51",
          7183 => x"56",
          7184 => x"83",
          7185 => x"39",
          7186 => x"19",
          7187 => x"83",
          7188 => x"0b",
          7189 => x"81",
          7190 => x"39",
          7191 => x"7c",
          7192 => x"74",
          7193 => x"38",
          7194 => x"7b",
          7195 => x"ec",
          7196 => x"08",
          7197 => x"06",
          7198 => x"81",
          7199 => x"8a",
          7200 => x"05",
          7201 => x"06",
          7202 => x"bf",
          7203 => x"38",
          7204 => x"55",
          7205 => x"7a",
          7206 => x"98",
          7207 => x"77",
          7208 => x"3f",
          7209 => x"08",
          7210 => x"98",
          7211 => x"82",
          7212 => x"81",
          7213 => x"38",
          7214 => x"ff",
          7215 => x"98",
          7216 => x"18",
          7217 => x"74",
          7218 => x"7e",
          7219 => x"08",
          7220 => x"2e",
          7221 => x"8d",
          7222 => x"ce",
          7223 => x"b6",
          7224 => x"ee",
          7225 => x"08",
          7226 => x"d1",
          7227 => x"b6",
          7228 => x"2e",
          7229 => x"82",
          7230 => x"1b",
          7231 => x"5a",
          7232 => x"2e",
          7233 => x"78",
          7234 => x"11",
          7235 => x"55",
          7236 => x"85",
          7237 => x"31",
          7238 => x"76",
          7239 => x"81",
          7240 => x"c8",
          7241 => x"b6",
          7242 => x"a6",
          7243 => x"11",
          7244 => x"56",
          7245 => x"27",
          7246 => x"80",
          7247 => x"08",
          7248 => x"2b",
          7249 => x"b4",
          7250 => x"b5",
          7251 => x"80",
          7252 => x"34",
          7253 => x"56",
          7254 => x"8c",
          7255 => x"19",
          7256 => x"38",
          7257 => x"b6",
          7258 => x"98",
          7259 => x"38",
          7260 => x"12",
          7261 => x"9c",
          7262 => x"18",
          7263 => x"06",
          7264 => x"31",
          7265 => x"76",
          7266 => x"7b",
          7267 => x"08",
          7268 => x"cd",
          7269 => x"b6",
          7270 => x"b6",
          7271 => x"7c",
          7272 => x"08",
          7273 => x"1f",
          7274 => x"cb",
          7275 => x"55",
          7276 => x"16",
          7277 => x"31",
          7278 => x"7f",
          7279 => x"94",
          7280 => x"70",
          7281 => x"8c",
          7282 => x"58",
          7283 => x"76",
          7284 => x"75",
          7285 => x"19",
          7286 => x"39",
          7287 => x"80",
          7288 => x"74",
          7289 => x"80",
          7290 => x"b6",
          7291 => x"3d",
          7292 => x"3d",
          7293 => x"3d",
          7294 => x"70",
          7295 => x"ea",
          7296 => x"98",
          7297 => x"b6",
          7298 => x"fb",
          7299 => x"33",
          7300 => x"70",
          7301 => x"55",
          7302 => x"2e",
          7303 => x"a0",
          7304 => x"78",
          7305 => x"3f",
          7306 => x"08",
          7307 => x"98",
          7308 => x"38",
          7309 => x"8b",
          7310 => x"07",
          7311 => x"8b",
          7312 => x"16",
          7313 => x"52",
          7314 => x"dd",
          7315 => x"16",
          7316 => x"15",
          7317 => x"3f",
          7318 => x"0a",
          7319 => x"51",
          7320 => x"76",
          7321 => x"51",
          7322 => x"78",
          7323 => x"83",
          7324 => x"51",
          7325 => x"82",
          7326 => x"90",
          7327 => x"bf",
          7328 => x"73",
          7329 => x"76",
          7330 => x"0c",
          7331 => x"04",
          7332 => x"76",
          7333 => x"fe",
          7334 => x"b6",
          7335 => x"82",
          7336 => x"9c",
          7337 => x"fc",
          7338 => x"51",
          7339 => x"82",
          7340 => x"53",
          7341 => x"08",
          7342 => x"b6",
          7343 => x"0c",
          7344 => x"98",
          7345 => x"0d",
          7346 => x"0d",
          7347 => x"e6",
          7348 => x"52",
          7349 => x"b6",
          7350 => x"8b",
          7351 => x"98",
          7352 => x"e4",
          7353 => x"71",
          7354 => x"0c",
          7355 => x"04",
          7356 => x"80",
          7357 => x"d0",
          7358 => x"3d",
          7359 => x"3f",
          7360 => x"08",
          7361 => x"98",
          7362 => x"38",
          7363 => x"52",
          7364 => x"05",
          7365 => x"3f",
          7366 => x"08",
          7367 => x"98",
          7368 => x"02",
          7369 => x"33",
          7370 => x"55",
          7371 => x"25",
          7372 => x"7a",
          7373 => x"54",
          7374 => x"a2",
          7375 => x"84",
          7376 => x"06",
          7377 => x"73",
          7378 => x"38",
          7379 => x"70",
          7380 => x"a8",
          7381 => x"98",
          7382 => x"0c",
          7383 => x"b6",
          7384 => x"2e",
          7385 => x"83",
          7386 => x"74",
          7387 => x"0c",
          7388 => x"04",
          7389 => x"6f",
          7390 => x"80",
          7391 => x"53",
          7392 => x"b8",
          7393 => x"3d",
          7394 => x"3f",
          7395 => x"08",
          7396 => x"98",
          7397 => x"38",
          7398 => x"7c",
          7399 => x"47",
          7400 => x"54",
          7401 => x"81",
          7402 => x"52",
          7403 => x"52",
          7404 => x"3f",
          7405 => x"08",
          7406 => x"98",
          7407 => x"38",
          7408 => x"51",
          7409 => x"82",
          7410 => x"57",
          7411 => x"08",
          7412 => x"69",
          7413 => x"da",
          7414 => x"b6",
          7415 => x"76",
          7416 => x"d5",
          7417 => x"b6",
          7418 => x"82",
          7419 => x"82",
          7420 => x"52",
          7421 => x"eb",
          7422 => x"98",
          7423 => x"b6",
          7424 => x"38",
          7425 => x"51",
          7426 => x"73",
          7427 => x"08",
          7428 => x"76",
          7429 => x"d6",
          7430 => x"b6",
          7431 => x"82",
          7432 => x"80",
          7433 => x"76",
          7434 => x"81",
          7435 => x"82",
          7436 => x"39",
          7437 => x"38",
          7438 => x"bc",
          7439 => x"51",
          7440 => x"76",
          7441 => x"11",
          7442 => x"51",
          7443 => x"73",
          7444 => x"38",
          7445 => x"55",
          7446 => x"16",
          7447 => x"56",
          7448 => x"38",
          7449 => x"73",
          7450 => x"90",
          7451 => x"2e",
          7452 => x"16",
          7453 => x"ff",
          7454 => x"ff",
          7455 => x"58",
          7456 => x"74",
          7457 => x"75",
          7458 => x"18",
          7459 => x"58",
          7460 => x"fe",
          7461 => x"7b",
          7462 => x"06",
          7463 => x"18",
          7464 => x"58",
          7465 => x"80",
          7466 => x"e4",
          7467 => x"29",
          7468 => x"05",
          7469 => x"33",
          7470 => x"56",
          7471 => x"2e",
          7472 => x"16",
          7473 => x"33",
          7474 => x"73",
          7475 => x"16",
          7476 => x"26",
          7477 => x"55",
          7478 => x"91",
          7479 => x"54",
          7480 => x"70",
          7481 => x"34",
          7482 => x"ec",
          7483 => x"70",
          7484 => x"34",
          7485 => x"09",
          7486 => x"38",
          7487 => x"39",
          7488 => x"19",
          7489 => x"33",
          7490 => x"05",
          7491 => x"78",
          7492 => x"80",
          7493 => x"82",
          7494 => x"9e",
          7495 => x"f7",
          7496 => x"7d",
          7497 => x"05",
          7498 => x"57",
          7499 => x"3f",
          7500 => x"08",
          7501 => x"98",
          7502 => x"38",
          7503 => x"53",
          7504 => x"38",
          7505 => x"54",
          7506 => x"92",
          7507 => x"33",
          7508 => x"70",
          7509 => x"54",
          7510 => x"38",
          7511 => x"15",
          7512 => x"70",
          7513 => x"58",
          7514 => x"82",
          7515 => x"8a",
          7516 => x"89",
          7517 => x"53",
          7518 => x"b7",
          7519 => x"ff",
          7520 => x"db",
          7521 => x"b6",
          7522 => x"15",
          7523 => x"53",
          7524 => x"db",
          7525 => x"b6",
          7526 => x"26",
          7527 => x"30",
          7528 => x"70",
          7529 => x"77",
          7530 => x"18",
          7531 => x"51",
          7532 => x"88",
          7533 => x"73",
          7534 => x"52",
          7535 => x"ca",
          7536 => x"98",
          7537 => x"b6",
          7538 => x"2e",
          7539 => x"82",
          7540 => x"ff",
          7541 => x"38",
          7542 => x"08",
          7543 => x"73",
          7544 => x"73",
          7545 => x"9c",
          7546 => x"27",
          7547 => x"75",
          7548 => x"16",
          7549 => x"17",
          7550 => x"33",
          7551 => x"70",
          7552 => x"55",
          7553 => x"80",
          7554 => x"73",
          7555 => x"cc",
          7556 => x"b6",
          7557 => x"82",
          7558 => x"94",
          7559 => x"98",
          7560 => x"39",
          7561 => x"51",
          7562 => x"82",
          7563 => x"54",
          7564 => x"be",
          7565 => x"27",
          7566 => x"53",
          7567 => x"08",
          7568 => x"73",
          7569 => x"ff",
          7570 => x"15",
          7571 => x"16",
          7572 => x"ff",
          7573 => x"80",
          7574 => x"73",
          7575 => x"c6",
          7576 => x"b6",
          7577 => x"38",
          7578 => x"16",
          7579 => x"80",
          7580 => x"0b",
          7581 => x"81",
          7582 => x"75",
          7583 => x"b6",
          7584 => x"58",
          7585 => x"54",
          7586 => x"74",
          7587 => x"73",
          7588 => x"90",
          7589 => x"c0",
          7590 => x"90",
          7591 => x"83",
          7592 => x"72",
          7593 => x"38",
          7594 => x"08",
          7595 => x"77",
          7596 => x"80",
          7597 => x"b6",
          7598 => x"3d",
          7599 => x"3d",
          7600 => x"89",
          7601 => x"2e",
          7602 => x"80",
          7603 => x"fc",
          7604 => x"3d",
          7605 => x"e1",
          7606 => x"b6",
          7607 => x"82",
          7608 => x"80",
          7609 => x"76",
          7610 => x"75",
          7611 => x"3f",
          7612 => x"08",
          7613 => x"98",
          7614 => x"38",
          7615 => x"70",
          7616 => x"57",
          7617 => x"a2",
          7618 => x"33",
          7619 => x"70",
          7620 => x"55",
          7621 => x"2e",
          7622 => x"16",
          7623 => x"51",
          7624 => x"82",
          7625 => x"88",
          7626 => x"54",
          7627 => x"84",
          7628 => x"52",
          7629 => x"e5",
          7630 => x"98",
          7631 => x"84",
          7632 => x"06",
          7633 => x"55",
          7634 => x"80",
          7635 => x"80",
          7636 => x"54",
          7637 => x"98",
          7638 => x"0d",
          7639 => x"0d",
          7640 => x"fc",
          7641 => x"52",
          7642 => x"3f",
          7643 => x"08",
          7644 => x"b6",
          7645 => x"0c",
          7646 => x"04",
          7647 => x"77",
          7648 => x"fc",
          7649 => x"53",
          7650 => x"de",
          7651 => x"98",
          7652 => x"b6",
          7653 => x"df",
          7654 => x"38",
          7655 => x"08",
          7656 => x"cd",
          7657 => x"b6",
          7658 => x"80",
          7659 => x"b6",
          7660 => x"73",
          7661 => x"3f",
          7662 => x"08",
          7663 => x"98",
          7664 => x"09",
          7665 => x"38",
          7666 => x"39",
          7667 => x"08",
          7668 => x"52",
          7669 => x"b3",
          7670 => x"73",
          7671 => x"3f",
          7672 => x"08",
          7673 => x"30",
          7674 => x"9f",
          7675 => x"b6",
          7676 => x"51",
          7677 => x"72",
          7678 => x"0c",
          7679 => x"04",
          7680 => x"65",
          7681 => x"89",
          7682 => x"96",
          7683 => x"df",
          7684 => x"b6",
          7685 => x"82",
          7686 => x"b2",
          7687 => x"75",
          7688 => x"3f",
          7689 => x"08",
          7690 => x"98",
          7691 => x"02",
          7692 => x"33",
          7693 => x"55",
          7694 => x"25",
          7695 => x"55",
          7696 => x"80",
          7697 => x"76",
          7698 => x"d4",
          7699 => x"82",
          7700 => x"94",
          7701 => x"f0",
          7702 => x"65",
          7703 => x"53",
          7704 => x"05",
          7705 => x"51",
          7706 => x"82",
          7707 => x"5b",
          7708 => x"08",
          7709 => x"7c",
          7710 => x"08",
          7711 => x"fe",
          7712 => x"08",
          7713 => x"55",
          7714 => x"91",
          7715 => x"0c",
          7716 => x"81",
          7717 => x"39",
          7718 => x"c7",
          7719 => x"98",
          7720 => x"55",
          7721 => x"2e",
          7722 => x"bf",
          7723 => x"5f",
          7724 => x"92",
          7725 => x"51",
          7726 => x"82",
          7727 => x"ff",
          7728 => x"82",
          7729 => x"81",
          7730 => x"82",
          7731 => x"30",
          7732 => x"98",
          7733 => x"25",
          7734 => x"19",
          7735 => x"5a",
          7736 => x"08",
          7737 => x"38",
          7738 => x"a4",
          7739 => x"b6",
          7740 => x"58",
          7741 => x"77",
          7742 => x"7d",
          7743 => x"bf",
          7744 => x"b6",
          7745 => x"82",
          7746 => x"80",
          7747 => x"70",
          7748 => x"ff",
          7749 => x"56",
          7750 => x"2e",
          7751 => x"9e",
          7752 => x"51",
          7753 => x"3f",
          7754 => x"08",
          7755 => x"06",
          7756 => x"80",
          7757 => x"19",
          7758 => x"54",
          7759 => x"14",
          7760 => x"c5",
          7761 => x"98",
          7762 => x"06",
          7763 => x"80",
          7764 => x"19",
          7765 => x"54",
          7766 => x"06",
          7767 => x"79",
          7768 => x"78",
          7769 => x"79",
          7770 => x"84",
          7771 => x"07",
          7772 => x"84",
          7773 => x"82",
          7774 => x"92",
          7775 => x"f9",
          7776 => x"8a",
          7777 => x"53",
          7778 => x"e3",
          7779 => x"b6",
          7780 => x"82",
          7781 => x"81",
          7782 => x"17",
          7783 => x"81",
          7784 => x"17",
          7785 => x"2a",
          7786 => x"51",
          7787 => x"55",
          7788 => x"81",
          7789 => x"17",
          7790 => x"8c",
          7791 => x"81",
          7792 => x"9b",
          7793 => x"98",
          7794 => x"17",
          7795 => x"51",
          7796 => x"82",
          7797 => x"74",
          7798 => x"56",
          7799 => x"98",
          7800 => x"76",
          7801 => x"c6",
          7802 => x"98",
          7803 => x"09",
          7804 => x"38",
          7805 => x"b6",
          7806 => x"2e",
          7807 => x"85",
          7808 => x"a3",
          7809 => x"38",
          7810 => x"b6",
          7811 => x"15",
          7812 => x"38",
          7813 => x"53",
          7814 => x"08",
          7815 => x"c3",
          7816 => x"b6",
          7817 => x"94",
          7818 => x"18",
          7819 => x"33",
          7820 => x"54",
          7821 => x"34",
          7822 => x"85",
          7823 => x"18",
          7824 => x"74",
          7825 => x"0c",
          7826 => x"04",
          7827 => x"82",
          7828 => x"ff",
          7829 => x"a1",
          7830 => x"e4",
          7831 => x"98",
          7832 => x"b6",
          7833 => x"f5",
          7834 => x"a1",
          7835 => x"95",
          7836 => x"58",
          7837 => x"82",
          7838 => x"55",
          7839 => x"08",
          7840 => x"02",
          7841 => x"33",
          7842 => x"70",
          7843 => x"55",
          7844 => x"73",
          7845 => x"75",
          7846 => x"80",
          7847 => x"bd",
          7848 => x"d6",
          7849 => x"81",
          7850 => x"87",
          7851 => x"ad",
          7852 => x"78",
          7853 => x"3f",
          7854 => x"08",
          7855 => x"70",
          7856 => x"55",
          7857 => x"2e",
          7858 => x"78",
          7859 => x"98",
          7860 => x"08",
          7861 => x"38",
          7862 => x"b6",
          7863 => x"76",
          7864 => x"70",
          7865 => x"b5",
          7866 => x"98",
          7867 => x"b6",
          7868 => x"e9",
          7869 => x"98",
          7870 => x"51",
          7871 => x"82",
          7872 => x"55",
          7873 => x"08",
          7874 => x"55",
          7875 => x"82",
          7876 => x"84",
          7877 => x"82",
          7878 => x"80",
          7879 => x"51",
          7880 => x"82",
          7881 => x"82",
          7882 => x"30",
          7883 => x"98",
          7884 => x"25",
          7885 => x"75",
          7886 => x"38",
          7887 => x"8f",
          7888 => x"75",
          7889 => x"c1",
          7890 => x"b6",
          7891 => x"74",
          7892 => x"51",
          7893 => x"3f",
          7894 => x"08",
          7895 => x"b6",
          7896 => x"3d",
          7897 => x"3d",
          7898 => x"99",
          7899 => x"52",
          7900 => x"d8",
          7901 => x"b6",
          7902 => x"82",
          7903 => x"82",
          7904 => x"5e",
          7905 => x"3d",
          7906 => x"cf",
          7907 => x"b6",
          7908 => x"82",
          7909 => x"86",
          7910 => x"82",
          7911 => x"b6",
          7912 => x"2e",
          7913 => x"82",
          7914 => x"80",
          7915 => x"70",
          7916 => x"06",
          7917 => x"54",
          7918 => x"38",
          7919 => x"52",
          7920 => x"52",
          7921 => x"3f",
          7922 => x"08",
          7923 => x"82",
          7924 => x"83",
          7925 => x"82",
          7926 => x"81",
          7927 => x"06",
          7928 => x"54",
          7929 => x"08",
          7930 => x"81",
          7931 => x"81",
          7932 => x"39",
          7933 => x"38",
          7934 => x"08",
          7935 => x"c4",
          7936 => x"b6",
          7937 => x"82",
          7938 => x"81",
          7939 => x"53",
          7940 => x"19",
          7941 => x"8c",
          7942 => x"ae",
          7943 => x"34",
          7944 => x"0b",
          7945 => x"82",
          7946 => x"52",
          7947 => x"51",
          7948 => x"3f",
          7949 => x"b4",
          7950 => x"c9",
          7951 => x"53",
          7952 => x"53",
          7953 => x"51",
          7954 => x"3f",
          7955 => x"0b",
          7956 => x"34",
          7957 => x"80",
          7958 => x"51",
          7959 => x"78",
          7960 => x"83",
          7961 => x"51",
          7962 => x"82",
          7963 => x"54",
          7964 => x"08",
          7965 => x"88",
          7966 => x"64",
          7967 => x"ff",
          7968 => x"75",
          7969 => x"78",
          7970 => x"3f",
          7971 => x"0b",
          7972 => x"78",
          7973 => x"83",
          7974 => x"51",
          7975 => x"3f",
          7976 => x"08",
          7977 => x"80",
          7978 => x"76",
          7979 => x"ae",
          7980 => x"b6",
          7981 => x"3d",
          7982 => x"3d",
          7983 => x"84",
          7984 => x"f1",
          7985 => x"a8",
          7986 => x"05",
          7987 => x"51",
          7988 => x"82",
          7989 => x"55",
          7990 => x"08",
          7991 => x"78",
          7992 => x"08",
          7993 => x"70",
          7994 => x"b8",
          7995 => x"98",
          7996 => x"b6",
          7997 => x"b9",
          7998 => x"9b",
          7999 => x"a0",
          8000 => x"55",
          8001 => x"38",
          8002 => x"3d",
          8003 => x"3d",
          8004 => x"51",
          8005 => x"3f",
          8006 => x"52",
          8007 => x"52",
          8008 => x"dd",
          8009 => x"08",
          8010 => x"cb",
          8011 => x"b6",
          8012 => x"82",
          8013 => x"95",
          8014 => x"2e",
          8015 => x"88",
          8016 => x"3d",
          8017 => x"38",
          8018 => x"e5",
          8019 => x"98",
          8020 => x"09",
          8021 => x"b8",
          8022 => x"c9",
          8023 => x"b6",
          8024 => x"82",
          8025 => x"81",
          8026 => x"56",
          8027 => x"3d",
          8028 => x"52",
          8029 => x"ff",
          8030 => x"02",
          8031 => x"8b",
          8032 => x"16",
          8033 => x"2a",
          8034 => x"51",
          8035 => x"89",
          8036 => x"07",
          8037 => x"17",
          8038 => x"81",
          8039 => x"34",
          8040 => x"70",
          8041 => x"81",
          8042 => x"55",
          8043 => x"80",
          8044 => x"64",
          8045 => x"38",
          8046 => x"51",
          8047 => x"82",
          8048 => x"52",
          8049 => x"b7",
          8050 => x"55",
          8051 => x"08",
          8052 => x"dd",
          8053 => x"98",
          8054 => x"51",
          8055 => x"3f",
          8056 => x"08",
          8057 => x"11",
          8058 => x"82",
          8059 => x"80",
          8060 => x"16",
          8061 => x"ae",
          8062 => x"06",
          8063 => x"53",
          8064 => x"51",
          8065 => x"78",
          8066 => x"83",
          8067 => x"39",
          8068 => x"08",
          8069 => x"51",
          8070 => x"82",
          8071 => x"55",
          8072 => x"08",
          8073 => x"51",
          8074 => x"3f",
          8075 => x"08",
          8076 => x"b6",
          8077 => x"3d",
          8078 => x"3d",
          8079 => x"db",
          8080 => x"84",
          8081 => x"05",
          8082 => x"82",
          8083 => x"d0",
          8084 => x"3d",
          8085 => x"3f",
          8086 => x"08",
          8087 => x"98",
          8088 => x"38",
          8089 => x"52",
          8090 => x"05",
          8091 => x"3f",
          8092 => x"08",
          8093 => x"98",
          8094 => x"02",
          8095 => x"33",
          8096 => x"54",
          8097 => x"aa",
          8098 => x"06",
          8099 => x"8b",
          8100 => x"06",
          8101 => x"07",
          8102 => x"56",
          8103 => x"34",
          8104 => x"0b",
          8105 => x"78",
          8106 => x"a9",
          8107 => x"98",
          8108 => x"82",
          8109 => x"95",
          8110 => x"ef",
          8111 => x"56",
          8112 => x"3d",
          8113 => x"94",
          8114 => x"f4",
          8115 => x"98",
          8116 => x"b6",
          8117 => x"cb",
          8118 => x"63",
          8119 => x"d4",
          8120 => x"c0",
          8121 => x"98",
          8122 => x"b6",
          8123 => x"38",
          8124 => x"05",
          8125 => x"06",
          8126 => x"73",
          8127 => x"16",
          8128 => x"22",
          8129 => x"07",
          8130 => x"1f",
          8131 => x"c2",
          8132 => x"81",
          8133 => x"34",
          8134 => x"b3",
          8135 => x"b6",
          8136 => x"74",
          8137 => x"0c",
          8138 => x"04",
          8139 => x"69",
          8140 => x"80",
          8141 => x"d0",
          8142 => x"3d",
          8143 => x"3f",
          8144 => x"08",
          8145 => x"08",
          8146 => x"b6",
          8147 => x"80",
          8148 => x"57",
          8149 => x"81",
          8150 => x"70",
          8151 => x"55",
          8152 => x"80",
          8153 => x"5d",
          8154 => x"52",
          8155 => x"52",
          8156 => x"a9",
          8157 => x"98",
          8158 => x"b6",
          8159 => x"d1",
          8160 => x"73",
          8161 => x"3f",
          8162 => x"08",
          8163 => x"98",
          8164 => x"82",
          8165 => x"82",
          8166 => x"65",
          8167 => x"78",
          8168 => x"7b",
          8169 => x"55",
          8170 => x"34",
          8171 => x"8a",
          8172 => x"38",
          8173 => x"1a",
          8174 => x"34",
          8175 => x"9e",
          8176 => x"70",
          8177 => x"51",
          8178 => x"a0",
          8179 => x"8e",
          8180 => x"2e",
          8181 => x"86",
          8182 => x"34",
          8183 => x"30",
          8184 => x"80",
          8185 => x"7a",
          8186 => x"c1",
          8187 => x"2e",
          8188 => x"a0",
          8189 => x"51",
          8190 => x"3f",
          8191 => x"08",
          8192 => x"98",
          8193 => x"7b",
          8194 => x"55",
          8195 => x"73",
          8196 => x"38",
          8197 => x"73",
          8198 => x"38",
          8199 => x"15",
          8200 => x"ff",
          8201 => x"82",
          8202 => x"7b",
          8203 => x"b6",
          8204 => x"3d",
          8205 => x"3d",
          8206 => x"9c",
          8207 => x"05",
          8208 => x"51",
          8209 => x"82",
          8210 => x"82",
          8211 => x"56",
          8212 => x"98",
          8213 => x"38",
          8214 => x"52",
          8215 => x"52",
          8216 => x"c0",
          8217 => x"70",
          8218 => x"ff",
          8219 => x"55",
          8220 => x"27",
          8221 => x"78",
          8222 => x"ff",
          8223 => x"05",
          8224 => x"55",
          8225 => x"3f",
          8226 => x"08",
          8227 => x"38",
          8228 => x"70",
          8229 => x"ff",
          8230 => x"82",
          8231 => x"80",
          8232 => x"74",
          8233 => x"07",
          8234 => x"4e",
          8235 => x"82",
          8236 => x"55",
          8237 => x"70",
          8238 => x"06",
          8239 => x"99",
          8240 => x"e0",
          8241 => x"ff",
          8242 => x"54",
          8243 => x"27",
          8244 => x"ae",
          8245 => x"55",
          8246 => x"a3",
          8247 => x"82",
          8248 => x"ff",
          8249 => x"82",
          8250 => x"93",
          8251 => x"75",
          8252 => x"76",
          8253 => x"38",
          8254 => x"77",
          8255 => x"86",
          8256 => x"39",
          8257 => x"27",
          8258 => x"88",
          8259 => x"78",
          8260 => x"5a",
          8261 => x"57",
          8262 => x"81",
          8263 => x"81",
          8264 => x"33",
          8265 => x"06",
          8266 => x"57",
          8267 => x"fe",
          8268 => x"3d",
          8269 => x"55",
          8270 => x"2e",
          8271 => x"76",
          8272 => x"38",
          8273 => x"55",
          8274 => x"33",
          8275 => x"a0",
          8276 => x"06",
          8277 => x"17",
          8278 => x"38",
          8279 => x"43",
          8280 => x"3d",
          8281 => x"ff",
          8282 => x"82",
          8283 => x"54",
          8284 => x"08",
          8285 => x"81",
          8286 => x"ff",
          8287 => x"82",
          8288 => x"54",
          8289 => x"08",
          8290 => x"80",
          8291 => x"54",
          8292 => x"80",
          8293 => x"b6",
          8294 => x"2e",
          8295 => x"80",
          8296 => x"54",
          8297 => x"80",
          8298 => x"52",
          8299 => x"bd",
          8300 => x"b6",
          8301 => x"82",
          8302 => x"b1",
          8303 => x"82",
          8304 => x"52",
          8305 => x"ab",
          8306 => x"54",
          8307 => x"15",
          8308 => x"78",
          8309 => x"ff",
          8310 => x"79",
          8311 => x"83",
          8312 => x"51",
          8313 => x"3f",
          8314 => x"08",
          8315 => x"74",
          8316 => x"0c",
          8317 => x"04",
          8318 => x"60",
          8319 => x"05",
          8320 => x"33",
          8321 => x"05",
          8322 => x"40",
          8323 => x"da",
          8324 => x"98",
          8325 => x"b6",
          8326 => x"bd",
          8327 => x"33",
          8328 => x"b5",
          8329 => x"2e",
          8330 => x"1a",
          8331 => x"90",
          8332 => x"33",
          8333 => x"70",
          8334 => x"55",
          8335 => x"38",
          8336 => x"97",
          8337 => x"82",
          8338 => x"58",
          8339 => x"7e",
          8340 => x"70",
          8341 => x"55",
          8342 => x"56",
          8343 => x"a4",
          8344 => x"7d",
          8345 => x"70",
          8346 => x"2a",
          8347 => x"08",
          8348 => x"08",
          8349 => x"5d",
          8350 => x"77",
          8351 => x"98",
          8352 => x"26",
          8353 => x"57",
          8354 => x"59",
          8355 => x"52",
          8356 => x"ae",
          8357 => x"15",
          8358 => x"98",
          8359 => x"26",
          8360 => x"55",
          8361 => x"08",
          8362 => x"99",
          8363 => x"98",
          8364 => x"ff",
          8365 => x"b6",
          8366 => x"38",
          8367 => x"75",
          8368 => x"81",
          8369 => x"93",
          8370 => x"80",
          8371 => x"2e",
          8372 => x"ff",
          8373 => x"58",
          8374 => x"7d",
          8375 => x"38",
          8376 => x"55",
          8377 => x"b4",
          8378 => x"56",
          8379 => x"09",
          8380 => x"38",
          8381 => x"53",
          8382 => x"51",
          8383 => x"3f",
          8384 => x"08",
          8385 => x"98",
          8386 => x"38",
          8387 => x"ff",
          8388 => x"5c",
          8389 => x"84",
          8390 => x"5c",
          8391 => x"12",
          8392 => x"80",
          8393 => x"78",
          8394 => x"7c",
          8395 => x"90",
          8396 => x"c0",
          8397 => x"90",
          8398 => x"15",
          8399 => x"90",
          8400 => x"54",
          8401 => x"91",
          8402 => x"31",
          8403 => x"84",
          8404 => x"07",
          8405 => x"16",
          8406 => x"73",
          8407 => x"0c",
          8408 => x"04",
          8409 => x"6b",
          8410 => x"05",
          8411 => x"33",
          8412 => x"5a",
          8413 => x"bd",
          8414 => x"80",
          8415 => x"98",
          8416 => x"f8",
          8417 => x"98",
          8418 => x"82",
          8419 => x"70",
          8420 => x"74",
          8421 => x"38",
          8422 => x"82",
          8423 => x"81",
          8424 => x"81",
          8425 => x"ff",
          8426 => x"82",
          8427 => x"81",
          8428 => x"81",
          8429 => x"83",
          8430 => x"c0",
          8431 => x"2a",
          8432 => x"51",
          8433 => x"74",
          8434 => x"99",
          8435 => x"53",
          8436 => x"51",
          8437 => x"3f",
          8438 => x"08",
          8439 => x"55",
          8440 => x"92",
          8441 => x"80",
          8442 => x"38",
          8443 => x"06",
          8444 => x"2e",
          8445 => x"48",
          8446 => x"87",
          8447 => x"79",
          8448 => x"78",
          8449 => x"26",
          8450 => x"19",
          8451 => x"74",
          8452 => x"38",
          8453 => x"e4",
          8454 => x"2a",
          8455 => x"70",
          8456 => x"59",
          8457 => x"7a",
          8458 => x"56",
          8459 => x"80",
          8460 => x"51",
          8461 => x"74",
          8462 => x"99",
          8463 => x"53",
          8464 => x"51",
          8465 => x"3f",
          8466 => x"b6",
          8467 => x"ac",
          8468 => x"2a",
          8469 => x"82",
          8470 => x"43",
          8471 => x"83",
          8472 => x"66",
          8473 => x"60",
          8474 => x"90",
          8475 => x"31",
          8476 => x"80",
          8477 => x"8a",
          8478 => x"56",
          8479 => x"26",
          8480 => x"77",
          8481 => x"81",
          8482 => x"74",
          8483 => x"38",
          8484 => x"55",
          8485 => x"83",
          8486 => x"81",
          8487 => x"80",
          8488 => x"38",
          8489 => x"55",
          8490 => x"5e",
          8491 => x"89",
          8492 => x"5a",
          8493 => x"09",
          8494 => x"e1",
          8495 => x"38",
          8496 => x"57",
          8497 => x"b1",
          8498 => x"5a",
          8499 => x"9d",
          8500 => x"26",
          8501 => x"b1",
          8502 => x"10",
          8503 => x"22",
          8504 => x"74",
          8505 => x"38",
          8506 => x"ee",
          8507 => x"66",
          8508 => x"90",
          8509 => x"98",
          8510 => x"84",
          8511 => x"89",
          8512 => x"a0",
          8513 => x"82",
          8514 => x"fc",
          8515 => x"56",
          8516 => x"f0",
          8517 => x"80",
          8518 => x"d3",
          8519 => x"38",
          8520 => x"57",
          8521 => x"b0",
          8522 => x"5a",
          8523 => x"9d",
          8524 => x"26",
          8525 => x"b0",
          8526 => x"10",
          8527 => x"22",
          8528 => x"74",
          8529 => x"38",
          8530 => x"ee",
          8531 => x"66",
          8532 => x"b0",
          8533 => x"98",
          8534 => x"05",
          8535 => x"98",
          8536 => x"26",
          8537 => x"0b",
          8538 => x"08",
          8539 => x"98",
          8540 => x"11",
          8541 => x"05",
          8542 => x"83",
          8543 => x"2a",
          8544 => x"a0",
          8545 => x"7d",
          8546 => x"69",
          8547 => x"05",
          8548 => x"72",
          8549 => x"5c",
          8550 => x"59",
          8551 => x"2e",
          8552 => x"89",
          8553 => x"60",
          8554 => x"84",
          8555 => x"5d",
          8556 => x"18",
          8557 => x"68",
          8558 => x"74",
          8559 => x"af",
          8560 => x"31",
          8561 => x"53",
          8562 => x"52",
          8563 => x"b4",
          8564 => x"98",
          8565 => x"83",
          8566 => x"06",
          8567 => x"b6",
          8568 => x"ff",
          8569 => x"dd",
          8570 => x"83",
          8571 => x"2a",
          8572 => x"be",
          8573 => x"39",
          8574 => x"09",
          8575 => x"c5",
          8576 => x"f5",
          8577 => x"98",
          8578 => x"38",
          8579 => x"79",
          8580 => x"80",
          8581 => x"38",
          8582 => x"96",
          8583 => x"06",
          8584 => x"2e",
          8585 => x"5e",
          8586 => x"82",
          8587 => x"9f",
          8588 => x"38",
          8589 => x"38",
          8590 => x"81",
          8591 => x"fc",
          8592 => x"ab",
          8593 => x"7d",
          8594 => x"81",
          8595 => x"7d",
          8596 => x"78",
          8597 => x"74",
          8598 => x"8e",
          8599 => x"9c",
          8600 => x"53",
          8601 => x"51",
          8602 => x"3f",
          8603 => x"af",
          8604 => x"51",
          8605 => x"3f",
          8606 => x"8b",
          8607 => x"a1",
          8608 => x"8d",
          8609 => x"83",
          8610 => x"52",
          8611 => x"ff",
          8612 => x"81",
          8613 => x"34",
          8614 => x"70",
          8615 => x"2a",
          8616 => x"54",
          8617 => x"1b",
          8618 => x"88",
          8619 => x"74",
          8620 => x"26",
          8621 => x"83",
          8622 => x"52",
          8623 => x"ff",
          8624 => x"8a",
          8625 => x"a0",
          8626 => x"a1",
          8627 => x"0b",
          8628 => x"bf",
          8629 => x"51",
          8630 => x"3f",
          8631 => x"9a",
          8632 => x"a0",
          8633 => x"52",
          8634 => x"ff",
          8635 => x"7d",
          8636 => x"81",
          8637 => x"38",
          8638 => x"0a",
          8639 => x"1b",
          8640 => x"ce",
          8641 => x"a4",
          8642 => x"a0",
          8643 => x"52",
          8644 => x"ff",
          8645 => x"81",
          8646 => x"51",
          8647 => x"3f",
          8648 => x"1b",
          8649 => x"8c",
          8650 => x"0b",
          8651 => x"34",
          8652 => x"c2",
          8653 => x"53",
          8654 => x"52",
          8655 => x"51",
          8656 => x"88",
          8657 => x"a7",
          8658 => x"a0",
          8659 => x"83",
          8660 => x"52",
          8661 => x"ff",
          8662 => x"ff",
          8663 => x"1c",
          8664 => x"a6",
          8665 => x"53",
          8666 => x"52",
          8667 => x"ff",
          8668 => x"82",
          8669 => x"83",
          8670 => x"52",
          8671 => x"b4",
          8672 => x"60",
          8673 => x"7e",
          8674 => x"d7",
          8675 => x"82",
          8676 => x"83",
          8677 => x"83",
          8678 => x"06",
          8679 => x"75",
          8680 => x"05",
          8681 => x"7e",
          8682 => x"b7",
          8683 => x"53",
          8684 => x"51",
          8685 => x"3f",
          8686 => x"a4",
          8687 => x"51",
          8688 => x"3f",
          8689 => x"e4",
          8690 => x"e4",
          8691 => x"9f",
          8692 => x"18",
          8693 => x"1b",
          8694 => x"f6",
          8695 => x"83",
          8696 => x"ff",
          8697 => x"82",
          8698 => x"78",
          8699 => x"c4",
          8700 => x"60",
          8701 => x"7a",
          8702 => x"ff",
          8703 => x"75",
          8704 => x"53",
          8705 => x"51",
          8706 => x"3f",
          8707 => x"52",
          8708 => x"9f",
          8709 => x"56",
          8710 => x"83",
          8711 => x"06",
          8712 => x"52",
          8713 => x"9e",
          8714 => x"52",
          8715 => x"ff",
          8716 => x"f0",
          8717 => x"1b",
          8718 => x"87",
          8719 => x"55",
          8720 => x"83",
          8721 => x"74",
          8722 => x"ff",
          8723 => x"7c",
          8724 => x"74",
          8725 => x"38",
          8726 => x"54",
          8727 => x"52",
          8728 => x"99",
          8729 => x"b6",
          8730 => x"87",
          8731 => x"53",
          8732 => x"08",
          8733 => x"ff",
          8734 => x"76",
          8735 => x"31",
          8736 => x"cd",
          8737 => x"58",
          8738 => x"ff",
          8739 => x"55",
          8740 => x"83",
          8741 => x"61",
          8742 => x"26",
          8743 => x"57",
          8744 => x"53",
          8745 => x"51",
          8746 => x"3f",
          8747 => x"08",
          8748 => x"76",
          8749 => x"31",
          8750 => x"db",
          8751 => x"7d",
          8752 => x"38",
          8753 => x"83",
          8754 => x"8a",
          8755 => x"7d",
          8756 => x"38",
          8757 => x"81",
          8758 => x"80",
          8759 => x"80",
          8760 => x"7a",
          8761 => x"bc",
          8762 => x"d5",
          8763 => x"ff",
          8764 => x"83",
          8765 => x"77",
          8766 => x"0b",
          8767 => x"81",
          8768 => x"34",
          8769 => x"34",
          8770 => x"34",
          8771 => x"56",
          8772 => x"52",
          8773 => x"b4",
          8774 => x"0b",
          8775 => x"82",
          8776 => x"82",
          8777 => x"56",
          8778 => x"34",
          8779 => x"08",
          8780 => x"60",
          8781 => x"1b",
          8782 => x"96",
          8783 => x"83",
          8784 => x"ff",
          8785 => x"81",
          8786 => x"7a",
          8787 => x"ff",
          8788 => x"81",
          8789 => x"98",
          8790 => x"80",
          8791 => x"7e",
          8792 => x"e3",
          8793 => x"82",
          8794 => x"90",
          8795 => x"8e",
          8796 => x"81",
          8797 => x"82",
          8798 => x"56",
          8799 => x"98",
          8800 => x"0d",
          8801 => x"0d",
          8802 => x"59",
          8803 => x"ff",
          8804 => x"57",
          8805 => x"b4",
          8806 => x"f8",
          8807 => x"81",
          8808 => x"52",
          8809 => x"dc",
          8810 => x"2e",
          8811 => x"9c",
          8812 => x"33",
          8813 => x"2e",
          8814 => x"76",
          8815 => x"58",
          8816 => x"57",
          8817 => x"09",
          8818 => x"38",
          8819 => x"78",
          8820 => x"38",
          8821 => x"82",
          8822 => x"8d",
          8823 => x"f7",
          8824 => x"02",
          8825 => x"05",
          8826 => x"77",
          8827 => x"81",
          8828 => x"8d",
          8829 => x"e7",
          8830 => x"08",
          8831 => x"24",
          8832 => x"17",
          8833 => x"8c",
          8834 => x"77",
          8835 => x"16",
          8836 => x"25",
          8837 => x"3d",
          8838 => x"75",
          8839 => x"52",
          8840 => x"cb",
          8841 => x"76",
          8842 => x"70",
          8843 => x"2a",
          8844 => x"51",
          8845 => x"84",
          8846 => x"19",
          8847 => x"8b",
          8848 => x"f9",
          8849 => x"84",
          8850 => x"56",
          8851 => x"a7",
          8852 => x"fc",
          8853 => x"53",
          8854 => x"75",
          8855 => x"a1",
          8856 => x"98",
          8857 => x"84",
          8858 => x"2e",
          8859 => x"87",
          8860 => x"08",
          8861 => x"ff",
          8862 => x"b6",
          8863 => x"3d",
          8864 => x"3d",
          8865 => x"80",
          8866 => x"52",
          8867 => x"9a",
          8868 => x"74",
          8869 => x"0d",
          8870 => x"0d",
          8871 => x"05",
          8872 => x"86",
          8873 => x"54",
          8874 => x"73",
          8875 => x"fe",
          8876 => x"51",
          8877 => x"98",
          8878 => x"00",
          8879 => x"ff",
          8880 => x"ff",
          8881 => x"00",
          8882 => x"ff",
          8883 => x"2b",
          8884 => x"2b",
          8885 => x"2b",
          8886 => x"2b",
          8887 => x"2b",
          8888 => x"2b",
          8889 => x"2b",
          8890 => x"2b",
          8891 => x"2b",
          8892 => x"2b",
          8893 => x"2b",
          8894 => x"2b",
          8895 => x"2b",
          8896 => x"2b",
          8897 => x"2b",
          8898 => x"2b",
          8899 => x"2b",
          8900 => x"2b",
          8901 => x"2b",
          8902 => x"2b",
          8903 => x"41",
          8904 => x"41",
          8905 => x"41",
          8906 => x"41",
          8907 => x"41",
          8908 => x"47",
          8909 => x"48",
          8910 => x"49",
          8911 => x"4b",
          8912 => x"48",
          8913 => x"46",
          8914 => x"4a",
          8915 => x"4b",
          8916 => x"4a",
          8917 => x"4b",
          8918 => x"4a",
          8919 => x"49",
          8920 => x"46",
          8921 => x"49",
          8922 => x"49",
          8923 => x"4a",
          8924 => x"46",
          8925 => x"46",
          8926 => x"4a",
          8927 => x"4b",
          8928 => x"4b",
          8929 => x"4b",
          8930 => x"0e",
          8931 => x"17",
          8932 => x"17",
          8933 => x"0e",
          8934 => x"17",
          8935 => x"17",
          8936 => x"17",
          8937 => x"17",
          8938 => x"17",
          8939 => x"17",
          8940 => x"17",
          8941 => x"0e",
          8942 => x"17",
          8943 => x"0e",
          8944 => x"0e",
          8945 => x"17",
          8946 => x"17",
          8947 => x"17",
          8948 => x"17",
          8949 => x"17",
          8950 => x"17",
          8951 => x"17",
          8952 => x"17",
          8953 => x"17",
          8954 => x"17",
          8955 => x"17",
          8956 => x"17",
          8957 => x"17",
          8958 => x"17",
          8959 => x"17",
          8960 => x"17",
          8961 => x"17",
          8962 => x"17",
          8963 => x"17",
          8964 => x"17",
          8965 => x"17",
          8966 => x"17",
          8967 => x"17",
          8968 => x"17",
          8969 => x"17",
          8970 => x"17",
          8971 => x"17",
          8972 => x"17",
          8973 => x"17",
          8974 => x"17",
          8975 => x"17",
          8976 => x"17",
          8977 => x"17",
          8978 => x"17",
          8979 => x"17",
          8980 => x"17",
          8981 => x"0f",
          8982 => x"17",
          8983 => x"17",
          8984 => x"17",
          8985 => x"17",
          8986 => x"11",
          8987 => x"17",
          8988 => x"17",
          8989 => x"17",
          8990 => x"17",
          8991 => x"17",
          8992 => x"17",
          8993 => x"17",
          8994 => x"17",
          8995 => x"17",
          8996 => x"17",
          8997 => x"0e",
          8998 => x"10",
          8999 => x"0e",
          9000 => x"0e",
          9001 => x"0e",
          9002 => x"17",
          9003 => x"10",
          9004 => x"17",
          9005 => x"17",
          9006 => x"0e",
          9007 => x"17",
          9008 => x"17",
          9009 => x"10",
          9010 => x"10",
          9011 => x"17",
          9012 => x"17",
          9013 => x"0f",
          9014 => x"17",
          9015 => x"11",
          9016 => x"17",
          9017 => x"17",
          9018 => x"11",
          9019 => x"6e",
          9020 => x"00",
          9021 => x"6f",
          9022 => x"00",
          9023 => x"6e",
          9024 => x"00",
          9025 => x"6f",
          9026 => x"00",
          9027 => x"78",
          9028 => x"00",
          9029 => x"6c",
          9030 => x"00",
          9031 => x"6f",
          9032 => x"00",
          9033 => x"69",
          9034 => x"00",
          9035 => x"75",
          9036 => x"00",
          9037 => x"62",
          9038 => x"68",
          9039 => x"77",
          9040 => x"64",
          9041 => x"65",
          9042 => x"64",
          9043 => x"65",
          9044 => x"6c",
          9045 => x"00",
          9046 => x"70",
          9047 => x"73",
          9048 => x"74",
          9049 => x"73",
          9050 => x"00",
          9051 => x"66",
          9052 => x"00",
          9053 => x"73",
          9054 => x"00",
          9055 => x"61",
          9056 => x"00",
          9057 => x"61",
          9058 => x"00",
          9059 => x"6c",
          9060 => x"00",
          9061 => x"00",
          9062 => x"73",
          9063 => x"72",
          9064 => x"00",
          9065 => x"74",
          9066 => x"61",
          9067 => x"72",
          9068 => x"2e",
          9069 => x"73",
          9070 => x"6f",
          9071 => x"65",
          9072 => x"2e",
          9073 => x"20",
          9074 => x"65",
          9075 => x"75",
          9076 => x"00",
          9077 => x"20",
          9078 => x"68",
          9079 => x"75",
          9080 => x"00",
          9081 => x"76",
          9082 => x"64",
          9083 => x"6c",
          9084 => x"6d",
          9085 => x"00",
          9086 => x"63",
          9087 => x"20",
          9088 => x"69",
          9089 => x"00",
          9090 => x"6c",
          9091 => x"6c",
          9092 => x"64",
          9093 => x"78",
          9094 => x"73",
          9095 => x"00",
          9096 => x"6c",
          9097 => x"61",
          9098 => x"65",
          9099 => x"76",
          9100 => x"64",
          9101 => x"00",
          9102 => x"20",
          9103 => x"77",
          9104 => x"65",
          9105 => x"6f",
          9106 => x"74",
          9107 => x"00",
          9108 => x"69",
          9109 => x"6e",
          9110 => x"65",
          9111 => x"73",
          9112 => x"76",
          9113 => x"64",
          9114 => x"00",
          9115 => x"73",
          9116 => x"6f",
          9117 => x"6e",
          9118 => x"65",
          9119 => x"00",
          9120 => x"20",
          9121 => x"70",
          9122 => x"62",
          9123 => x"66",
          9124 => x"73",
          9125 => x"65",
          9126 => x"6f",
          9127 => x"20",
          9128 => x"64",
          9129 => x"2e",
          9130 => x"72",
          9131 => x"20",
          9132 => x"72",
          9133 => x"2e",
          9134 => x"6d",
          9135 => x"74",
          9136 => x"70",
          9137 => x"74",
          9138 => x"20",
          9139 => x"63",
          9140 => x"65",
          9141 => x"00",
          9142 => x"6c",
          9143 => x"73",
          9144 => x"63",
          9145 => x"2e",
          9146 => x"73",
          9147 => x"69",
          9148 => x"6e",
          9149 => x"65",
          9150 => x"79",
          9151 => x"00",
          9152 => x"6f",
          9153 => x"6e",
          9154 => x"70",
          9155 => x"66",
          9156 => x"73",
          9157 => x"00",
          9158 => x"72",
          9159 => x"74",
          9160 => x"20",
          9161 => x"6f",
          9162 => x"63",
          9163 => x"00",
          9164 => x"63",
          9165 => x"73",
          9166 => x"00",
          9167 => x"6b",
          9168 => x"6e",
          9169 => x"72",
          9170 => x"00",
          9171 => x"6c",
          9172 => x"79",
          9173 => x"20",
          9174 => x"61",
          9175 => x"6c",
          9176 => x"79",
          9177 => x"2f",
          9178 => x"2e",
          9179 => x"00",
          9180 => x"61",
          9181 => x"00",
          9182 => x"25",
          9183 => x"78",
          9184 => x"3d",
          9185 => x"6c",
          9186 => x"32",
          9187 => x"38",
          9188 => x"20",
          9189 => x"42",
          9190 => x"38",
          9191 => x"25",
          9192 => x"78",
          9193 => x"38",
          9194 => x"00",
          9195 => x"38",
          9196 => x"00",
          9197 => x"20",
          9198 => x"34",
          9199 => x"00",
          9200 => x"20",
          9201 => x"20",
          9202 => x"00",
          9203 => x"32",
          9204 => x"00",
          9205 => x"00",
          9206 => x"00",
          9207 => x"00",
          9208 => x"53",
          9209 => x"2a",
          9210 => x"20",
          9211 => x"00",
          9212 => x"2f",
          9213 => x"32",
          9214 => x"00",
          9215 => x"2e",
          9216 => x"00",
          9217 => x"50",
          9218 => x"72",
          9219 => x"25",
          9220 => x"29",
          9221 => x"20",
          9222 => x"2a",
          9223 => x"00",
          9224 => x"55",
          9225 => x"74",
          9226 => x"75",
          9227 => x"48",
          9228 => x"6c",
          9229 => x"00",
          9230 => x"6d",
          9231 => x"69",
          9232 => x"72",
          9233 => x"74",
          9234 => x"32",
          9235 => x"74",
          9236 => x"75",
          9237 => x"00",
          9238 => x"43",
          9239 => x"52",
          9240 => x"6e",
          9241 => x"72",
          9242 => x"00",
          9243 => x"43",
          9244 => x"57",
          9245 => x"6e",
          9246 => x"72",
          9247 => x"00",
          9248 => x"52",
          9249 => x"52",
          9250 => x"6e",
          9251 => x"72",
          9252 => x"00",
          9253 => x"52",
          9254 => x"54",
          9255 => x"6e",
          9256 => x"72",
          9257 => x"00",
          9258 => x"52",
          9259 => x"52",
          9260 => x"6e",
          9261 => x"72",
          9262 => x"00",
          9263 => x"52",
          9264 => x"54",
          9265 => x"6e",
          9266 => x"72",
          9267 => x"00",
          9268 => x"74",
          9269 => x"67",
          9270 => x"20",
          9271 => x"65",
          9272 => x"2e",
          9273 => x"61",
          9274 => x"6e",
          9275 => x"69",
          9276 => x"2e",
          9277 => x"00",
          9278 => x"74",
          9279 => x"65",
          9280 => x"61",
          9281 => x"00",
          9282 => x"53",
          9283 => x"74",
          9284 => x"00",
          9285 => x"69",
          9286 => x"20",
          9287 => x"69",
          9288 => x"69",
          9289 => x"73",
          9290 => x"64",
          9291 => x"72",
          9292 => x"2c",
          9293 => x"65",
          9294 => x"20",
          9295 => x"74",
          9296 => x"6e",
          9297 => x"6c",
          9298 => x"00",
          9299 => x"00",
          9300 => x"65",
          9301 => x"6e",
          9302 => x"2e",
          9303 => x"00",
          9304 => x"70",
          9305 => x"67",
          9306 => x"00",
          9307 => x"6d",
          9308 => x"69",
          9309 => x"2e",
          9310 => x"00",
          9311 => x"38",
          9312 => x"25",
          9313 => x"29",
          9314 => x"30",
          9315 => x"28",
          9316 => x"78",
          9317 => x"00",
          9318 => x"6d",
          9319 => x"65",
          9320 => x"79",
          9321 => x"6f",
          9322 => x"65",
          9323 => x"00",
          9324 => x"38",
          9325 => x"25",
          9326 => x"2d",
          9327 => x"3f",
          9328 => x"38",
          9329 => x"25",
          9330 => x"2d",
          9331 => x"38",
          9332 => x"25",
          9333 => x"58",
          9334 => x"00",
          9335 => x"65",
          9336 => x"69",
          9337 => x"63",
          9338 => x"20",
          9339 => x"30",
          9340 => x"20",
          9341 => x"0a",
          9342 => x"6c",
          9343 => x"67",
          9344 => x"64",
          9345 => x"20",
          9346 => x"6c",
          9347 => x"2e",
          9348 => x"00",
          9349 => x"6c",
          9350 => x"65",
          9351 => x"6e",
          9352 => x"63",
          9353 => x"20",
          9354 => x"29",
          9355 => x"00",
          9356 => x"73",
          9357 => x"74",
          9358 => x"20",
          9359 => x"6c",
          9360 => x"74",
          9361 => x"2e",
          9362 => x"00",
          9363 => x"6c",
          9364 => x"65",
          9365 => x"74",
          9366 => x"2e",
          9367 => x"00",
          9368 => x"55",
          9369 => x"6e",
          9370 => x"3a",
          9371 => x"5c",
          9372 => x"25",
          9373 => x"00",
          9374 => x"3a",
          9375 => x"5c",
          9376 => x"00",
          9377 => x"3a",
          9378 => x"00",
          9379 => x"64",
          9380 => x"6d",
          9381 => x"64",
          9382 => x"00",
          9383 => x"6e",
          9384 => x"67",
          9385 => x"00",
          9386 => x"61",
          9387 => x"6e",
          9388 => x"6e",
          9389 => x"72",
          9390 => x"73",
          9391 => x"00",
          9392 => x"2f",
          9393 => x"25",
          9394 => x"64",
          9395 => x"3a",
          9396 => x"25",
          9397 => x"0a",
          9398 => x"43",
          9399 => x"6e",
          9400 => x"75",
          9401 => x"69",
          9402 => x"00",
          9403 => x"66",
          9404 => x"20",
          9405 => x"20",
          9406 => x"66",
          9407 => x"00",
          9408 => x"44",
          9409 => x"63",
          9410 => x"69",
          9411 => x"65",
          9412 => x"74",
          9413 => x"00",
          9414 => x"20",
          9415 => x"20",
          9416 => x"41",
          9417 => x"28",
          9418 => x"58",
          9419 => x"38",
          9420 => x"0a",
          9421 => x"20",
          9422 => x"52",
          9423 => x"20",
          9424 => x"28",
          9425 => x"58",
          9426 => x"38",
          9427 => x"0a",
          9428 => x"20",
          9429 => x"53",
          9430 => x"52",
          9431 => x"28",
          9432 => x"58",
          9433 => x"38",
          9434 => x"0a",
          9435 => x"20",
          9436 => x"41",
          9437 => x"20",
          9438 => x"28",
          9439 => x"58",
          9440 => x"38",
          9441 => x"0a",
          9442 => x"20",
          9443 => x"4d",
          9444 => x"20",
          9445 => x"28",
          9446 => x"58",
          9447 => x"38",
          9448 => x"0a",
          9449 => x"20",
          9450 => x"20",
          9451 => x"44",
          9452 => x"28",
          9453 => x"69",
          9454 => x"20",
          9455 => x"32",
          9456 => x"0a",
          9457 => x"20",
          9458 => x"4d",
          9459 => x"20",
          9460 => x"28",
          9461 => x"65",
          9462 => x"20",
          9463 => x"32",
          9464 => x"0a",
          9465 => x"20",
          9466 => x"54",
          9467 => x"54",
          9468 => x"28",
          9469 => x"6e",
          9470 => x"73",
          9471 => x"32",
          9472 => x"0a",
          9473 => x"20",
          9474 => x"53",
          9475 => x"4e",
          9476 => x"55",
          9477 => x"00",
          9478 => x"20",
          9479 => x"20",
          9480 => x"00",
          9481 => x"20",
          9482 => x"43",
          9483 => x"00",
          9484 => x"20",
          9485 => x"32",
          9486 => x"20",
          9487 => x"49",
          9488 => x"64",
          9489 => x"73",
          9490 => x"00",
          9491 => x"20",
          9492 => x"55",
          9493 => x"73",
          9494 => x"56",
          9495 => x"6f",
          9496 => x"64",
          9497 => x"73",
          9498 => x"20",
          9499 => x"58",
          9500 => x"00",
          9501 => x"20",
          9502 => x"55",
          9503 => x"6d",
          9504 => x"20",
          9505 => x"72",
          9506 => x"64",
          9507 => x"73",
          9508 => x"20",
          9509 => x"58",
          9510 => x"00",
          9511 => x"20",
          9512 => x"61",
          9513 => x"53",
          9514 => x"74",
          9515 => x"64",
          9516 => x"73",
          9517 => x"20",
          9518 => x"20",
          9519 => x"58",
          9520 => x"00",
          9521 => x"73",
          9522 => x"00",
          9523 => x"20",
          9524 => x"55",
          9525 => x"20",
          9526 => x"20",
          9527 => x"20",
          9528 => x"20",
          9529 => x"20",
          9530 => x"20",
          9531 => x"58",
          9532 => x"00",
          9533 => x"20",
          9534 => x"73",
          9535 => x"20",
          9536 => x"63",
          9537 => x"72",
          9538 => x"20",
          9539 => x"20",
          9540 => x"20",
          9541 => x"25",
          9542 => x"4d",
          9543 => x"00",
          9544 => x"20",
          9545 => x"52",
          9546 => x"43",
          9547 => x"6b",
          9548 => x"65",
          9549 => x"20",
          9550 => x"20",
          9551 => x"20",
          9552 => x"25",
          9553 => x"4d",
          9554 => x"00",
          9555 => x"20",
          9556 => x"73",
          9557 => x"6e",
          9558 => x"44",
          9559 => x"20",
          9560 => x"63",
          9561 => x"72",
          9562 => x"20",
          9563 => x"25",
          9564 => x"4d",
          9565 => x"00",
          9566 => x"61",
          9567 => x"00",
          9568 => x"64",
          9569 => x"00",
          9570 => x"65",
          9571 => x"00",
          9572 => x"4f",
          9573 => x"4f",
          9574 => x"00",
          9575 => x"6b",
          9576 => x"6e",
          9577 => x"97",
          9578 => x"00",
          9579 => x"00",
          9580 => x"96",
          9581 => x"00",
          9582 => x"00",
          9583 => x"96",
          9584 => x"00",
          9585 => x"00",
          9586 => x"96",
          9587 => x"00",
          9588 => x"00",
          9589 => x"96",
          9590 => x"00",
          9591 => x"00",
          9592 => x"96",
          9593 => x"00",
          9594 => x"00",
          9595 => x"96",
          9596 => x"00",
          9597 => x"00",
          9598 => x"96",
          9599 => x"00",
          9600 => x"00",
          9601 => x"96",
          9602 => x"00",
          9603 => x"00",
          9604 => x"96",
          9605 => x"00",
          9606 => x"00",
          9607 => x"96",
          9608 => x"00",
          9609 => x"00",
          9610 => x"96",
          9611 => x"00",
          9612 => x"00",
          9613 => x"96",
          9614 => x"00",
          9615 => x"00",
          9616 => x"96",
          9617 => x"00",
          9618 => x"00",
          9619 => x"96",
          9620 => x"00",
          9621 => x"00",
          9622 => x"96",
          9623 => x"00",
          9624 => x"00",
          9625 => x"96",
          9626 => x"00",
          9627 => x"00",
          9628 => x"96",
          9629 => x"00",
          9630 => x"00",
          9631 => x"96",
          9632 => x"00",
          9633 => x"00",
          9634 => x"96",
          9635 => x"00",
          9636 => x"00",
          9637 => x"96",
          9638 => x"00",
          9639 => x"00",
          9640 => x"96",
          9641 => x"00",
          9642 => x"00",
          9643 => x"44",
          9644 => x"43",
          9645 => x"42",
          9646 => x"41",
          9647 => x"36",
          9648 => x"35",
          9649 => x"34",
          9650 => x"46",
          9651 => x"33",
          9652 => x"32",
          9653 => x"31",
          9654 => x"00",
          9655 => x"00",
          9656 => x"00",
          9657 => x"00",
          9658 => x"00",
          9659 => x"00",
          9660 => x"00",
          9661 => x"00",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"73",
          9666 => x"79",
          9667 => x"73",
          9668 => x"00",
          9669 => x"00",
          9670 => x"34",
          9671 => x"20",
          9672 => x"00",
          9673 => x"69",
          9674 => x"20",
          9675 => x"72",
          9676 => x"74",
          9677 => x"65",
          9678 => x"73",
          9679 => x"79",
          9680 => x"6c",
          9681 => x"6f",
          9682 => x"46",
          9683 => x"00",
          9684 => x"6e",
          9685 => x"20",
          9686 => x"6e",
          9687 => x"65",
          9688 => x"20",
          9689 => x"74",
          9690 => x"20",
          9691 => x"65",
          9692 => x"69",
          9693 => x"6c",
          9694 => x"2e",
          9695 => x"00",
          9696 => x"2b",
          9697 => x"3c",
          9698 => x"5b",
          9699 => x"00",
          9700 => x"54",
          9701 => x"54",
          9702 => x"00",
          9703 => x"90",
          9704 => x"4f",
          9705 => x"30",
          9706 => x"20",
          9707 => x"45",
          9708 => x"20",
          9709 => x"33",
          9710 => x"20",
          9711 => x"20",
          9712 => x"45",
          9713 => x"20",
          9714 => x"20",
          9715 => x"20",
          9716 => x"97",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"45",
          9721 => x"8f",
          9722 => x"45",
          9723 => x"8e",
          9724 => x"92",
          9725 => x"55",
          9726 => x"9a",
          9727 => x"9e",
          9728 => x"4f",
          9729 => x"a6",
          9730 => x"aa",
          9731 => x"ae",
          9732 => x"b2",
          9733 => x"b6",
          9734 => x"ba",
          9735 => x"be",
          9736 => x"c2",
          9737 => x"c6",
          9738 => x"ca",
          9739 => x"ce",
          9740 => x"d2",
          9741 => x"d6",
          9742 => x"da",
          9743 => x"de",
          9744 => x"e2",
          9745 => x"e6",
          9746 => x"ea",
          9747 => x"ee",
          9748 => x"f2",
          9749 => x"f6",
          9750 => x"fa",
          9751 => x"fe",
          9752 => x"2c",
          9753 => x"5d",
          9754 => x"2a",
          9755 => x"3f",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"02",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"8c",
          9767 => x"01",
          9768 => x"00",
          9769 => x"00",
          9770 => x"8c",
          9771 => x"01",
          9772 => x"00",
          9773 => x"00",
          9774 => x"8c",
          9775 => x"03",
          9776 => x"00",
          9777 => x"00",
          9778 => x"8d",
          9779 => x"03",
          9780 => x"00",
          9781 => x"00",
          9782 => x"8d",
          9783 => x"03",
          9784 => x"00",
          9785 => x"00",
          9786 => x"8d",
          9787 => x"04",
          9788 => x"00",
          9789 => x"00",
          9790 => x"8d",
          9791 => x"04",
          9792 => x"00",
          9793 => x"00",
          9794 => x"8d",
          9795 => x"04",
          9796 => x"00",
          9797 => x"00",
          9798 => x"8d",
          9799 => x"04",
          9800 => x"00",
          9801 => x"00",
          9802 => x"8d",
          9803 => x"04",
          9804 => x"00",
          9805 => x"00",
          9806 => x"8d",
          9807 => x"04",
          9808 => x"00",
          9809 => x"00",
          9810 => x"8d",
          9811 => x"04",
          9812 => x"00",
          9813 => x"00",
          9814 => x"8d",
          9815 => x"05",
          9816 => x"00",
          9817 => x"00",
          9818 => x"8d",
          9819 => x"05",
          9820 => x"00",
          9821 => x"00",
          9822 => x"8d",
          9823 => x"05",
          9824 => x"00",
          9825 => x"00",
          9826 => x"8d",
          9827 => x"05",
          9828 => x"00",
          9829 => x"00",
          9830 => x"8d",
          9831 => x"07",
          9832 => x"00",
          9833 => x"00",
          9834 => x"8d",
          9835 => x"07",
          9836 => x"00",
          9837 => x"00",
          9838 => x"8d",
          9839 => x"08",
          9840 => x"00",
          9841 => x"00",
          9842 => x"8d",
          9843 => x"08",
          9844 => x"00",
          9845 => x"00",
          9846 => x"8d",
          9847 => x"08",
          9848 => x"00",
          9849 => x"00",
          9850 => x"8d",
          9851 => x"08",
          9852 => x"00",
          9853 => x"00",
          9854 => x"8d",
          9855 => x"09",
          9856 => x"00",
          9857 => x"00",
          9858 => x"8d",
          9859 => x"09",
          9860 => x"00",
          9861 => x"00",
          9862 => x"8d",
          9863 => x"09",
          9864 => x"00",
          9865 => x"00",
          9866 => x"8d",
          9867 => x"09",
          9868 => x"00",
          9869 => x"00",
          9870 => x"00",
          9871 => x"00",
          9872 => x"7f",
          9873 => x"00",
          9874 => x"7f",
          9875 => x"00",
          9876 => x"7f",
          9877 => x"00",
          9878 => x"00",
          9879 => x"00",
          9880 => x"ff",
          9881 => x"00",
          9882 => x"00",
          9883 => x"78",
          9884 => x"00",
          9885 => x"e1",
          9886 => x"e1",
          9887 => x"e1",
          9888 => x"00",
          9889 => x"01",
          9890 => x"01",
          9891 => x"10",
          9892 => x"00",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"00",
          9898 => x"00",
          9899 => x"00",
          9900 => x"00",
          9901 => x"00",
          9902 => x"00",
          9903 => x"00",
          9904 => x"00",
          9905 => x"00",
          9906 => x"00",
          9907 => x"00",
          9908 => x"00",
          9909 => x"00",
          9910 => x"00",
          9911 => x"00",
          9912 => x"00",
          9913 => x"00",
          9914 => x"00",
          9915 => x"00",
          9916 => x"00",
          9917 => x"97",
          9918 => x"00",
          9919 => x"97",
          9920 => x"00",
          9921 => x"97",
          9922 => x"00",
          9923 => x"00",
          9924 => x"00",
          9925 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"85",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"82",
           389 => x"82",
           390 => x"b3",
           391 => x"b6",
           392 => x"d0",
           393 => x"b6",
           394 => x"e3",
           395 => x"a4",
           396 => x"90",
           397 => x"a4",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"82",
           403 => x"82",
           404 => x"82",
           405 => x"b1",
           406 => x"b6",
           407 => x"d0",
           408 => x"b6",
           409 => x"cf",
           410 => x"b6",
           411 => x"d0",
           412 => x"b6",
           413 => x"c9",
           414 => x"b6",
           415 => x"d0",
           416 => x"b6",
           417 => x"d8",
           418 => x"a4",
           419 => x"90",
           420 => x"a4",
           421 => x"2d",
           422 => x"08",
           423 => x"04",
           424 => x"0c",
           425 => x"82",
           426 => x"82",
           427 => x"82",
           428 => x"80",
           429 => x"82",
           430 => x"82",
           431 => x"82",
           432 => x"80",
           433 => x"82",
           434 => x"82",
           435 => x"82",
           436 => x"80",
           437 => x"82",
           438 => x"82",
           439 => x"82",
           440 => x"80",
           441 => x"82",
           442 => x"82",
           443 => x"82",
           444 => x"80",
           445 => x"82",
           446 => x"82",
           447 => x"82",
           448 => x"81",
           449 => x"82",
           450 => x"82",
           451 => x"82",
           452 => x"81",
           453 => x"82",
           454 => x"82",
           455 => x"82",
           456 => x"81",
           457 => x"82",
           458 => x"82",
           459 => x"82",
           460 => x"81",
           461 => x"82",
           462 => x"82",
           463 => x"82",
           464 => x"81",
           465 => x"82",
           466 => x"82",
           467 => x"82",
           468 => x"81",
           469 => x"82",
           470 => x"82",
           471 => x"82",
           472 => x"81",
           473 => x"82",
           474 => x"82",
           475 => x"82",
           476 => x"81",
           477 => x"82",
           478 => x"82",
           479 => x"82",
           480 => x"81",
           481 => x"82",
           482 => x"82",
           483 => x"82",
           484 => x"81",
           485 => x"82",
           486 => x"82",
           487 => x"82",
           488 => x"81",
           489 => x"82",
           490 => x"82",
           491 => x"82",
           492 => x"81",
           493 => x"82",
           494 => x"82",
           495 => x"82",
           496 => x"81",
           497 => x"82",
           498 => x"82",
           499 => x"82",
           500 => x"81",
           501 => x"82",
           502 => x"82",
           503 => x"82",
           504 => x"81",
           505 => x"82",
           506 => x"82",
           507 => x"82",
           508 => x"81",
           509 => x"82",
           510 => x"82",
           511 => x"82",
           512 => x"81",
           513 => x"82",
           514 => x"82",
           515 => x"82",
           516 => x"81",
           517 => x"82",
           518 => x"82",
           519 => x"82",
           520 => x"81",
           521 => x"82",
           522 => x"82",
           523 => x"82",
           524 => x"81",
           525 => x"82",
           526 => x"82",
           527 => x"82",
           528 => x"81",
           529 => x"82",
           530 => x"82",
           531 => x"82",
           532 => x"82",
           533 => x"82",
           534 => x"82",
           535 => x"82",
           536 => x"82",
           537 => x"82",
           538 => x"82",
           539 => x"82",
           540 => x"81",
           541 => x"82",
           542 => x"82",
           543 => x"82",
           544 => x"82",
           545 => x"82",
           546 => x"82",
           547 => x"82",
           548 => x"82",
           549 => x"82",
           550 => x"82",
           551 => x"82",
           552 => x"82",
           553 => x"82",
           554 => x"82",
           555 => x"82",
           556 => x"81",
           557 => x"82",
           558 => x"82",
           559 => x"82",
           560 => x"81",
           561 => x"82",
           562 => x"82",
           563 => x"82",
           564 => x"81",
           565 => x"82",
           566 => x"82",
           567 => x"82",
           568 => x"80",
           569 => x"82",
           570 => x"82",
           571 => x"82",
           572 => x"80",
           573 => x"82",
           574 => x"82",
           575 => x"82",
           576 => x"80",
           577 => x"82",
           578 => x"82",
           579 => x"82",
           580 => x"80",
           581 => x"82",
           582 => x"82",
           583 => x"82",
           584 => x"81",
           585 => x"82",
           586 => x"82",
           587 => x"82",
           588 => x"81",
           589 => x"82",
           590 => x"82",
           591 => x"82",
           592 => x"81",
           593 => x"82",
           594 => x"82",
           595 => x"82",
           596 => x"81",
           597 => x"82",
           598 => x"82",
           599 => x"3c",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"51",
           609 => x"73",
           610 => x"73",
           611 => x"81",
           612 => x"10",
           613 => x"07",
           614 => x"0c",
           615 => x"72",
           616 => x"81",
           617 => x"09",
           618 => x"71",
           619 => x"0a",
           620 => x"72",
           621 => x"51",
           622 => x"82",
           623 => x"82",
           624 => x"8e",
           625 => x"70",
           626 => x"0c",
           627 => x"93",
           628 => x"81",
           629 => x"86",
           630 => x"b6",
           631 => x"82",
           632 => x"fb",
           633 => x"b6",
           634 => x"05",
           635 => x"a4",
           636 => x"0c",
           637 => x"08",
           638 => x"54",
           639 => x"08",
           640 => x"53",
           641 => x"08",
           642 => x"9a",
           643 => x"98",
           644 => x"b6",
           645 => x"05",
           646 => x"a4",
           647 => x"08",
           648 => x"98",
           649 => x"87",
           650 => x"b6",
           651 => x"82",
           652 => x"02",
           653 => x"0c",
           654 => x"82",
           655 => x"90",
           656 => x"11",
           657 => x"32",
           658 => x"51",
           659 => x"71",
           660 => x"0b",
           661 => x"08",
           662 => x"25",
           663 => x"39",
           664 => x"b6",
           665 => x"05",
           666 => x"39",
           667 => x"08",
           668 => x"ff",
           669 => x"a4",
           670 => x"0c",
           671 => x"b6",
           672 => x"05",
           673 => x"a4",
           674 => x"08",
           675 => x"08",
           676 => x"82",
           677 => x"f8",
           678 => x"2e",
           679 => x"80",
           680 => x"a4",
           681 => x"08",
           682 => x"38",
           683 => x"08",
           684 => x"51",
           685 => x"82",
           686 => x"70",
           687 => x"08",
           688 => x"52",
           689 => x"08",
           690 => x"ff",
           691 => x"06",
           692 => x"0b",
           693 => x"08",
           694 => x"80",
           695 => x"b6",
           696 => x"05",
           697 => x"a4",
           698 => x"08",
           699 => x"73",
           700 => x"a4",
           701 => x"08",
           702 => x"b6",
           703 => x"05",
           704 => x"a4",
           705 => x"08",
           706 => x"b6",
           707 => x"05",
           708 => x"39",
           709 => x"08",
           710 => x"52",
           711 => x"82",
           712 => x"88",
           713 => x"82",
           714 => x"f4",
           715 => x"82",
           716 => x"f4",
           717 => x"b6",
           718 => x"3d",
           719 => x"a4",
           720 => x"b6",
           721 => x"82",
           722 => x"f4",
           723 => x"0b",
           724 => x"08",
           725 => x"82",
           726 => x"88",
           727 => x"b6",
           728 => x"05",
           729 => x"0b",
           730 => x"08",
           731 => x"82",
           732 => x"90",
           733 => x"b6",
           734 => x"05",
           735 => x"a4",
           736 => x"08",
           737 => x"a4",
           738 => x"08",
           739 => x"a4",
           740 => x"70",
           741 => x"81",
           742 => x"b6",
           743 => x"82",
           744 => x"dc",
           745 => x"b6",
           746 => x"05",
           747 => x"a4",
           748 => x"08",
           749 => x"80",
           750 => x"b6",
           751 => x"05",
           752 => x"b6",
           753 => x"8e",
           754 => x"b6",
           755 => x"82",
           756 => x"02",
           757 => x"0c",
           758 => x"82",
           759 => x"90",
           760 => x"b6",
           761 => x"05",
           762 => x"a4",
           763 => x"08",
           764 => x"a4",
           765 => x"08",
           766 => x"a4",
           767 => x"08",
           768 => x"3f",
           769 => x"08",
           770 => x"a4",
           771 => x"0c",
           772 => x"08",
           773 => x"70",
           774 => x"0c",
           775 => x"3d",
           776 => x"a4",
           777 => x"b6",
           778 => x"82",
           779 => x"ed",
           780 => x"0b",
           781 => x"08",
           782 => x"82",
           783 => x"88",
           784 => x"80",
           785 => x"0c",
           786 => x"08",
           787 => x"85",
           788 => x"81",
           789 => x"32",
           790 => x"51",
           791 => x"53",
           792 => x"8d",
           793 => x"82",
           794 => x"e0",
           795 => x"ac",
           796 => x"a4",
           797 => x"08",
           798 => x"53",
           799 => x"a4",
           800 => x"34",
           801 => x"06",
           802 => x"2e",
           803 => x"82",
           804 => x"8c",
           805 => x"05",
           806 => x"08",
           807 => x"82",
           808 => x"e4",
           809 => x"81",
           810 => x"72",
           811 => x"8b",
           812 => x"a4",
           813 => x"33",
           814 => x"27",
           815 => x"82",
           816 => x"f8",
           817 => x"72",
           818 => x"ee",
           819 => x"a4",
           820 => x"33",
           821 => x"2e",
           822 => x"80",
           823 => x"b6",
           824 => x"05",
           825 => x"2b",
           826 => x"51",
           827 => x"b2",
           828 => x"a4",
           829 => x"22",
           830 => x"70",
           831 => x"81",
           832 => x"51",
           833 => x"2e",
           834 => x"b6",
           835 => x"05",
           836 => x"80",
           837 => x"72",
           838 => x"08",
           839 => x"fe",
           840 => x"b6",
           841 => x"05",
           842 => x"2b",
           843 => x"70",
           844 => x"72",
           845 => x"51",
           846 => x"51",
           847 => x"82",
           848 => x"e8",
           849 => x"b6",
           850 => x"05",
           851 => x"b6",
           852 => x"05",
           853 => x"d0",
           854 => x"53",
           855 => x"a4",
           856 => x"34",
           857 => x"08",
           858 => x"70",
           859 => x"98",
           860 => x"53",
           861 => x"8b",
           862 => x"0b",
           863 => x"08",
           864 => x"82",
           865 => x"e4",
           866 => x"83",
           867 => x"06",
           868 => x"72",
           869 => x"82",
           870 => x"e8",
           871 => x"88",
           872 => x"2b",
           873 => x"70",
           874 => x"51",
           875 => x"72",
           876 => x"08",
           877 => x"fd",
           878 => x"b6",
           879 => x"05",
           880 => x"2a",
           881 => x"51",
           882 => x"80",
           883 => x"82",
           884 => x"e8",
           885 => x"98",
           886 => x"2c",
           887 => x"72",
           888 => x"0b",
           889 => x"08",
           890 => x"82",
           891 => x"f8",
           892 => x"11",
           893 => x"08",
           894 => x"53",
           895 => x"08",
           896 => x"80",
           897 => x"94",
           898 => x"a4",
           899 => x"08",
           900 => x"82",
           901 => x"70",
           902 => x"51",
           903 => x"82",
           904 => x"e4",
           905 => x"90",
           906 => x"72",
           907 => x"08",
           908 => x"82",
           909 => x"e4",
           910 => x"a0",
           911 => x"72",
           912 => x"08",
           913 => x"fc",
           914 => x"b6",
           915 => x"05",
           916 => x"80",
           917 => x"72",
           918 => x"08",
           919 => x"fc",
           920 => x"b6",
           921 => x"05",
           922 => x"c0",
           923 => x"72",
           924 => x"08",
           925 => x"fb",
           926 => x"b6",
           927 => x"05",
           928 => x"07",
           929 => x"82",
           930 => x"e4",
           931 => x"0b",
           932 => x"08",
           933 => x"fb",
           934 => x"b6",
           935 => x"05",
           936 => x"07",
           937 => x"82",
           938 => x"e4",
           939 => x"c1",
           940 => x"82",
           941 => x"fc",
           942 => x"b6",
           943 => x"05",
           944 => x"51",
           945 => x"b6",
           946 => x"05",
           947 => x"0b",
           948 => x"08",
           949 => x"8d",
           950 => x"b6",
           951 => x"05",
           952 => x"a4",
           953 => x"08",
           954 => x"b6",
           955 => x"05",
           956 => x"51",
           957 => x"b6",
           958 => x"05",
           959 => x"a4",
           960 => x"22",
           961 => x"53",
           962 => x"a4",
           963 => x"23",
           964 => x"82",
           965 => x"90",
           966 => x"b6",
           967 => x"05",
           968 => x"82",
           969 => x"90",
           970 => x"08",
           971 => x"08",
           972 => x"82",
           973 => x"e4",
           974 => x"83",
           975 => x"06",
           976 => x"53",
           977 => x"ab",
           978 => x"a4",
           979 => x"33",
           980 => x"53",
           981 => x"53",
           982 => x"08",
           983 => x"52",
           984 => x"3f",
           985 => x"08",
           986 => x"b6",
           987 => x"05",
           988 => x"82",
           989 => x"fc",
           990 => x"9d",
           991 => x"b6",
           992 => x"72",
           993 => x"08",
           994 => x"82",
           995 => x"ec",
           996 => x"82",
           997 => x"f4",
           998 => x"71",
           999 => x"72",
          1000 => x"08",
          1001 => x"8b",
          1002 => x"b6",
          1003 => x"05",
          1004 => x"a4",
          1005 => x"08",
          1006 => x"b6",
          1007 => x"05",
          1008 => x"82",
          1009 => x"fc",
          1010 => x"b6",
          1011 => x"05",
          1012 => x"2a",
          1013 => x"51",
          1014 => x"72",
          1015 => x"38",
          1016 => x"08",
          1017 => x"70",
          1018 => x"72",
          1019 => x"82",
          1020 => x"fc",
          1021 => x"53",
          1022 => x"82",
          1023 => x"53",
          1024 => x"a4",
          1025 => x"23",
          1026 => x"b6",
          1027 => x"05",
          1028 => x"f3",
          1029 => x"98",
          1030 => x"82",
          1031 => x"f4",
          1032 => x"b6",
          1033 => x"05",
          1034 => x"b6",
          1035 => x"05",
          1036 => x"31",
          1037 => x"82",
          1038 => x"ec",
          1039 => x"c1",
          1040 => x"a4",
          1041 => x"22",
          1042 => x"70",
          1043 => x"51",
          1044 => x"2e",
          1045 => x"b6",
          1046 => x"05",
          1047 => x"a4",
          1048 => x"08",
          1049 => x"b6",
          1050 => x"05",
          1051 => x"82",
          1052 => x"dc",
          1053 => x"a2",
          1054 => x"a4",
          1055 => x"08",
          1056 => x"08",
          1057 => x"84",
          1058 => x"a4",
          1059 => x"0c",
          1060 => x"b6",
          1061 => x"05",
          1062 => x"b6",
          1063 => x"05",
          1064 => x"a4",
          1065 => x"0c",
          1066 => x"08",
          1067 => x"80",
          1068 => x"82",
          1069 => x"e4",
          1070 => x"82",
          1071 => x"72",
          1072 => x"08",
          1073 => x"82",
          1074 => x"fc",
          1075 => x"82",
          1076 => x"fc",
          1077 => x"b6",
          1078 => x"05",
          1079 => x"bf",
          1080 => x"72",
          1081 => x"08",
          1082 => x"81",
          1083 => x"0b",
          1084 => x"08",
          1085 => x"a9",
          1086 => x"a4",
          1087 => x"22",
          1088 => x"07",
          1089 => x"82",
          1090 => x"e4",
          1091 => x"f8",
          1092 => x"a4",
          1093 => x"34",
          1094 => x"b6",
          1095 => x"05",
          1096 => x"a4",
          1097 => x"22",
          1098 => x"70",
          1099 => x"51",
          1100 => x"2e",
          1101 => x"b6",
          1102 => x"05",
          1103 => x"a4",
          1104 => x"08",
          1105 => x"b6",
          1106 => x"05",
          1107 => x"82",
          1108 => x"d8",
          1109 => x"a2",
          1110 => x"a4",
          1111 => x"08",
          1112 => x"08",
          1113 => x"84",
          1114 => x"a4",
          1115 => x"0c",
          1116 => x"b6",
          1117 => x"05",
          1118 => x"b6",
          1119 => x"05",
          1120 => x"a4",
          1121 => x"0c",
          1122 => x"08",
          1123 => x"70",
          1124 => x"53",
          1125 => x"a4",
          1126 => x"23",
          1127 => x"0b",
          1128 => x"08",
          1129 => x"82",
          1130 => x"f0",
          1131 => x"b6",
          1132 => x"05",
          1133 => x"a4",
          1134 => x"08",
          1135 => x"54",
          1136 => x"a3",
          1137 => x"b6",
          1138 => x"72",
          1139 => x"b6",
          1140 => x"05",
          1141 => x"a4",
          1142 => x"0c",
          1143 => x"08",
          1144 => x"70",
          1145 => x"89",
          1146 => x"38",
          1147 => x"08",
          1148 => x"53",
          1149 => x"82",
          1150 => x"f8",
          1151 => x"15",
          1152 => x"51",
          1153 => x"b6",
          1154 => x"05",
          1155 => x"82",
          1156 => x"f0",
          1157 => x"72",
          1158 => x"51",
          1159 => x"b6",
          1160 => x"05",
          1161 => x"a4",
          1162 => x"08",
          1163 => x"a4",
          1164 => x"33",
          1165 => x"b6",
          1166 => x"05",
          1167 => x"82",
          1168 => x"f0",
          1169 => x"b6",
          1170 => x"05",
          1171 => x"82",
          1172 => x"fc",
          1173 => x"53",
          1174 => x"82",
          1175 => x"70",
          1176 => x"08",
          1177 => x"53",
          1178 => x"08",
          1179 => x"80",
          1180 => x"fe",
          1181 => x"b6",
          1182 => x"05",
          1183 => x"a8",
          1184 => x"54",
          1185 => x"31",
          1186 => x"82",
          1187 => x"fc",
          1188 => x"b6",
          1189 => x"05",
          1190 => x"06",
          1191 => x"80",
          1192 => x"82",
          1193 => x"ec",
          1194 => x"11",
          1195 => x"82",
          1196 => x"ec",
          1197 => x"b6",
          1198 => x"05",
          1199 => x"2a",
          1200 => x"51",
          1201 => x"80",
          1202 => x"38",
          1203 => x"08",
          1204 => x"70",
          1205 => x"b6",
          1206 => x"05",
          1207 => x"a4",
          1208 => x"08",
          1209 => x"b6",
          1210 => x"05",
          1211 => x"a4",
          1212 => x"22",
          1213 => x"90",
          1214 => x"06",
          1215 => x"b6",
          1216 => x"05",
          1217 => x"53",
          1218 => x"a4",
          1219 => x"23",
          1220 => x"b6",
          1221 => x"05",
          1222 => x"53",
          1223 => x"a4",
          1224 => x"23",
          1225 => x"08",
          1226 => x"82",
          1227 => x"ec",
          1228 => x"b6",
          1229 => x"05",
          1230 => x"2a",
          1231 => x"51",
          1232 => x"80",
          1233 => x"38",
          1234 => x"08",
          1235 => x"70",
          1236 => x"98",
          1237 => x"a4",
          1238 => x"33",
          1239 => x"53",
          1240 => x"97",
          1241 => x"a4",
          1242 => x"22",
          1243 => x"51",
          1244 => x"b6",
          1245 => x"05",
          1246 => x"82",
          1247 => x"e8",
          1248 => x"82",
          1249 => x"fc",
          1250 => x"71",
          1251 => x"72",
          1252 => x"08",
          1253 => x"82",
          1254 => x"e4",
          1255 => x"83",
          1256 => x"06",
          1257 => x"72",
          1258 => x"38",
          1259 => x"08",
          1260 => x"70",
          1261 => x"90",
          1262 => x"2c",
          1263 => x"51",
          1264 => x"53",
          1265 => x"b6",
          1266 => x"05",
          1267 => x"31",
          1268 => x"82",
          1269 => x"ec",
          1270 => x"39",
          1271 => x"08",
          1272 => x"70",
          1273 => x"90",
          1274 => x"2c",
          1275 => x"51",
          1276 => x"53",
          1277 => x"b6",
          1278 => x"05",
          1279 => x"31",
          1280 => x"82",
          1281 => x"ec",
          1282 => x"b6",
          1283 => x"05",
          1284 => x"80",
          1285 => x"72",
          1286 => x"b6",
          1287 => x"05",
          1288 => x"54",
          1289 => x"b6",
          1290 => x"05",
          1291 => x"2b",
          1292 => x"51",
          1293 => x"25",
          1294 => x"b6",
          1295 => x"05",
          1296 => x"51",
          1297 => x"d2",
          1298 => x"a4",
          1299 => x"22",
          1300 => x"70",
          1301 => x"51",
          1302 => x"2e",
          1303 => x"b6",
          1304 => x"05",
          1305 => x"51",
          1306 => x"80",
          1307 => x"b6",
          1308 => x"05",
          1309 => x"2a",
          1310 => x"51",
          1311 => x"80",
          1312 => x"82",
          1313 => x"88",
          1314 => x"ab",
          1315 => x"3f",
          1316 => x"b6",
          1317 => x"05",
          1318 => x"2a",
          1319 => x"51",
          1320 => x"80",
          1321 => x"82",
          1322 => x"88",
          1323 => x"a0",
          1324 => x"3f",
          1325 => x"08",
          1326 => x"70",
          1327 => x"81",
          1328 => x"53",
          1329 => x"b1",
          1330 => x"a4",
          1331 => x"08",
          1332 => x"89",
          1333 => x"b6",
          1334 => x"05",
          1335 => x"90",
          1336 => x"06",
          1337 => x"b6",
          1338 => x"05",
          1339 => x"b6",
          1340 => x"05",
          1341 => x"bc",
          1342 => x"a4",
          1343 => x"22",
          1344 => x"70",
          1345 => x"51",
          1346 => x"2e",
          1347 => x"b6",
          1348 => x"05",
          1349 => x"54",
          1350 => x"b6",
          1351 => x"05",
          1352 => x"2b",
          1353 => x"51",
          1354 => x"25",
          1355 => x"b6",
          1356 => x"05",
          1357 => x"51",
          1358 => x"d2",
          1359 => x"a4",
          1360 => x"22",
          1361 => x"70",
          1362 => x"51",
          1363 => x"2e",
          1364 => x"b6",
          1365 => x"05",
          1366 => x"54",
          1367 => x"b6",
          1368 => x"05",
          1369 => x"2b",
          1370 => x"51",
          1371 => x"25",
          1372 => x"b6",
          1373 => x"05",
          1374 => x"51",
          1375 => x"d2",
          1376 => x"a4",
          1377 => x"22",
          1378 => x"70",
          1379 => x"51",
          1380 => x"38",
          1381 => x"08",
          1382 => x"ff",
          1383 => x"72",
          1384 => x"08",
          1385 => x"73",
          1386 => x"90",
          1387 => x"80",
          1388 => x"38",
          1389 => x"08",
          1390 => x"52",
          1391 => x"f4",
          1392 => x"82",
          1393 => x"f8",
          1394 => x"72",
          1395 => x"09",
          1396 => x"38",
          1397 => x"08",
          1398 => x"52",
          1399 => x"08",
          1400 => x"51",
          1401 => x"81",
          1402 => x"b6",
          1403 => x"05",
          1404 => x"80",
          1405 => x"81",
          1406 => x"38",
          1407 => x"08",
          1408 => x"ff",
          1409 => x"72",
          1410 => x"08",
          1411 => x"72",
          1412 => x"06",
          1413 => x"ff",
          1414 => x"bb",
          1415 => x"a4",
          1416 => x"08",
          1417 => x"a4",
          1418 => x"08",
          1419 => x"82",
          1420 => x"fc",
          1421 => x"05",
          1422 => x"08",
          1423 => x"53",
          1424 => x"ff",
          1425 => x"b6",
          1426 => x"05",
          1427 => x"80",
          1428 => x"81",
          1429 => x"38",
          1430 => x"08",
          1431 => x"ff",
          1432 => x"72",
          1433 => x"08",
          1434 => x"72",
          1435 => x"06",
          1436 => x"ff",
          1437 => x"df",
          1438 => x"a4",
          1439 => x"08",
          1440 => x"a4",
          1441 => x"08",
          1442 => x"53",
          1443 => x"82",
          1444 => x"fc",
          1445 => x"05",
          1446 => x"08",
          1447 => x"ff",
          1448 => x"b6",
          1449 => x"05",
          1450 => x"a8",
          1451 => x"82",
          1452 => x"88",
          1453 => x"82",
          1454 => x"f0",
          1455 => x"05",
          1456 => x"08",
          1457 => x"82",
          1458 => x"f0",
          1459 => x"33",
          1460 => x"e0",
          1461 => x"82",
          1462 => x"e4",
          1463 => x"87",
          1464 => x"06",
          1465 => x"72",
          1466 => x"c3",
          1467 => x"a4",
          1468 => x"22",
          1469 => x"54",
          1470 => x"a4",
          1471 => x"23",
          1472 => x"70",
          1473 => x"53",
          1474 => x"a3",
          1475 => x"a4",
          1476 => x"08",
          1477 => x"85",
          1478 => x"39",
          1479 => x"08",
          1480 => x"52",
          1481 => x"08",
          1482 => x"51",
          1483 => x"80",
          1484 => x"a4",
          1485 => x"23",
          1486 => x"82",
          1487 => x"f8",
          1488 => x"72",
          1489 => x"81",
          1490 => x"81",
          1491 => x"a4",
          1492 => x"23",
          1493 => x"b6",
          1494 => x"05",
          1495 => x"82",
          1496 => x"e8",
          1497 => x"0b",
          1498 => x"08",
          1499 => x"ea",
          1500 => x"b6",
          1501 => x"05",
          1502 => x"b6",
          1503 => x"05",
          1504 => x"b0",
          1505 => x"39",
          1506 => x"08",
          1507 => x"8c",
          1508 => x"82",
          1509 => x"e0",
          1510 => x"53",
          1511 => x"08",
          1512 => x"82",
          1513 => x"95",
          1514 => x"b6",
          1515 => x"82",
          1516 => x"02",
          1517 => x"0c",
          1518 => x"82",
          1519 => x"53",
          1520 => x"08",
          1521 => x"52",
          1522 => x"08",
          1523 => x"51",
          1524 => x"82",
          1525 => x"70",
          1526 => x"0c",
          1527 => x"0d",
          1528 => x"0c",
          1529 => x"a4",
          1530 => x"b6",
          1531 => x"3d",
          1532 => x"82",
          1533 => x"f8",
          1534 => x"cd",
          1535 => x"11",
          1536 => x"2a",
          1537 => x"70",
          1538 => x"51",
          1539 => x"72",
          1540 => x"38",
          1541 => x"b6",
          1542 => x"05",
          1543 => x"39",
          1544 => x"08",
          1545 => x"53",
          1546 => x"b6",
          1547 => x"05",
          1548 => x"82",
          1549 => x"88",
          1550 => x"72",
          1551 => x"08",
          1552 => x"72",
          1553 => x"53",
          1554 => x"b0",
          1555 => x"ec",
          1556 => x"ec",
          1557 => x"b6",
          1558 => x"05",
          1559 => x"11",
          1560 => x"72",
          1561 => x"98",
          1562 => x"80",
          1563 => x"38",
          1564 => x"b6",
          1565 => x"05",
          1566 => x"39",
          1567 => x"08",
          1568 => x"08",
          1569 => x"51",
          1570 => x"53",
          1571 => x"b6",
          1572 => x"72",
          1573 => x"38",
          1574 => x"b6",
          1575 => x"05",
          1576 => x"a4",
          1577 => x"08",
          1578 => x"a4",
          1579 => x"0c",
          1580 => x"a4",
          1581 => x"08",
          1582 => x"0c",
          1583 => x"82",
          1584 => x"04",
          1585 => x"08",
          1586 => x"a4",
          1587 => x"0d",
          1588 => x"b6",
          1589 => x"05",
          1590 => x"a4",
          1591 => x"08",
          1592 => x"70",
          1593 => x"81",
          1594 => x"06",
          1595 => x"51",
          1596 => x"2e",
          1597 => x"0b",
          1598 => x"08",
          1599 => x"80",
          1600 => x"b6",
          1601 => x"05",
          1602 => x"33",
          1603 => x"08",
          1604 => x"81",
          1605 => x"a4",
          1606 => x"0c",
          1607 => x"b6",
          1608 => x"05",
          1609 => x"ff",
          1610 => x"80",
          1611 => x"82",
          1612 => x"8c",
          1613 => x"b6",
          1614 => x"05",
          1615 => x"b6",
          1616 => x"05",
          1617 => x"11",
          1618 => x"72",
          1619 => x"98",
          1620 => x"80",
          1621 => x"38",
          1622 => x"b6",
          1623 => x"05",
          1624 => x"39",
          1625 => x"08",
          1626 => x"70",
          1627 => x"08",
          1628 => x"53",
          1629 => x"08",
          1630 => x"82",
          1631 => x"87",
          1632 => x"b6",
          1633 => x"82",
          1634 => x"02",
          1635 => x"0c",
          1636 => x"82",
          1637 => x"52",
          1638 => x"08",
          1639 => x"51",
          1640 => x"b6",
          1641 => x"82",
          1642 => x"53",
          1643 => x"82",
          1644 => x"04",
          1645 => x"08",
          1646 => x"a4",
          1647 => x"0d",
          1648 => x"08",
          1649 => x"85",
          1650 => x"81",
          1651 => x"32",
          1652 => x"51",
          1653 => x"53",
          1654 => x"8d",
          1655 => x"82",
          1656 => x"fc",
          1657 => x"cb",
          1658 => x"a4",
          1659 => x"08",
          1660 => x"70",
          1661 => x"81",
          1662 => x"51",
          1663 => x"2e",
          1664 => x"82",
          1665 => x"8c",
          1666 => x"b6",
          1667 => x"05",
          1668 => x"8c",
          1669 => x"14",
          1670 => x"38",
          1671 => x"08",
          1672 => x"70",
          1673 => x"b6",
          1674 => x"05",
          1675 => x"54",
          1676 => x"34",
          1677 => x"05",
          1678 => x"b6",
          1679 => x"05",
          1680 => x"08",
          1681 => x"12",
          1682 => x"a4",
          1683 => x"08",
          1684 => x"a4",
          1685 => x"0c",
          1686 => x"d7",
          1687 => x"a4",
          1688 => x"08",
          1689 => x"08",
          1690 => x"53",
          1691 => x"08",
          1692 => x"70",
          1693 => x"53",
          1694 => x"51",
          1695 => x"2d",
          1696 => x"08",
          1697 => x"38",
          1698 => x"08",
          1699 => x"8c",
          1700 => x"05",
          1701 => x"82",
          1702 => x"88",
          1703 => x"82",
          1704 => x"fc",
          1705 => x"53",
          1706 => x"0b",
          1707 => x"08",
          1708 => x"82",
          1709 => x"fc",
          1710 => x"b6",
          1711 => x"3d",
          1712 => x"a4",
          1713 => x"b6",
          1714 => x"82",
          1715 => x"f9",
          1716 => x"b6",
          1717 => x"05",
          1718 => x"33",
          1719 => x"70",
          1720 => x"51",
          1721 => x"80",
          1722 => x"ff",
          1723 => x"a4",
          1724 => x"0c",
          1725 => x"82",
          1726 => x"88",
          1727 => x"11",
          1728 => x"2a",
          1729 => x"51",
          1730 => x"71",
          1731 => x"c5",
          1732 => x"a4",
          1733 => x"08",
          1734 => x"08",
          1735 => x"53",
          1736 => x"33",
          1737 => x"06",
          1738 => x"85",
          1739 => x"b6",
          1740 => x"05",
          1741 => x"08",
          1742 => x"12",
          1743 => x"a4",
          1744 => x"08",
          1745 => x"70",
          1746 => x"08",
          1747 => x"51",
          1748 => x"b6",
          1749 => x"a4",
          1750 => x"08",
          1751 => x"70",
          1752 => x"81",
          1753 => x"51",
          1754 => x"2e",
          1755 => x"82",
          1756 => x"88",
          1757 => x"08",
          1758 => x"b6",
          1759 => x"05",
          1760 => x"82",
          1761 => x"fc",
          1762 => x"38",
          1763 => x"08",
          1764 => x"82",
          1765 => x"88",
          1766 => x"53",
          1767 => x"70",
          1768 => x"52",
          1769 => x"34",
          1770 => x"b6",
          1771 => x"05",
          1772 => x"39",
          1773 => x"08",
          1774 => x"70",
          1775 => x"71",
          1776 => x"a1",
          1777 => x"a4",
          1778 => x"08",
          1779 => x"08",
          1780 => x"52",
          1781 => x"51",
          1782 => x"82",
          1783 => x"70",
          1784 => x"08",
          1785 => x"52",
          1786 => x"08",
          1787 => x"80",
          1788 => x"38",
          1789 => x"08",
          1790 => x"82",
          1791 => x"f4",
          1792 => x"b6",
          1793 => x"05",
          1794 => x"33",
          1795 => x"08",
          1796 => x"52",
          1797 => x"08",
          1798 => x"ff",
          1799 => x"06",
          1800 => x"b6",
          1801 => x"05",
          1802 => x"52",
          1803 => x"a4",
          1804 => x"34",
          1805 => x"b6",
          1806 => x"05",
          1807 => x"52",
          1808 => x"a4",
          1809 => x"34",
          1810 => x"08",
          1811 => x"52",
          1812 => x"08",
          1813 => x"85",
          1814 => x"0b",
          1815 => x"08",
          1816 => x"a6",
          1817 => x"a4",
          1818 => x"08",
          1819 => x"81",
          1820 => x"0c",
          1821 => x"08",
          1822 => x"70",
          1823 => x"70",
          1824 => x"08",
          1825 => x"51",
          1826 => x"b6",
          1827 => x"05",
          1828 => x"98",
          1829 => x"0d",
          1830 => x"0c",
          1831 => x"a4",
          1832 => x"b6",
          1833 => x"3d",
          1834 => x"a4",
          1835 => x"08",
          1836 => x"08",
          1837 => x"82",
          1838 => x"8c",
          1839 => x"b6",
          1840 => x"05",
          1841 => x"a4",
          1842 => x"08",
          1843 => x"a2",
          1844 => x"a4",
          1845 => x"08",
          1846 => x"08",
          1847 => x"26",
          1848 => x"82",
          1849 => x"f8",
          1850 => x"b6",
          1851 => x"05",
          1852 => x"82",
          1853 => x"fc",
          1854 => x"27",
          1855 => x"82",
          1856 => x"fc",
          1857 => x"b6",
          1858 => x"05",
          1859 => x"b6",
          1860 => x"05",
          1861 => x"a4",
          1862 => x"08",
          1863 => x"08",
          1864 => x"05",
          1865 => x"08",
          1866 => x"82",
          1867 => x"90",
          1868 => x"05",
          1869 => x"08",
          1870 => x"82",
          1871 => x"90",
          1872 => x"05",
          1873 => x"08",
          1874 => x"82",
          1875 => x"90",
          1876 => x"2e",
          1877 => x"82",
          1878 => x"fc",
          1879 => x"05",
          1880 => x"08",
          1881 => x"82",
          1882 => x"f8",
          1883 => x"05",
          1884 => x"08",
          1885 => x"82",
          1886 => x"fc",
          1887 => x"b6",
          1888 => x"05",
          1889 => x"71",
          1890 => x"ff",
          1891 => x"b6",
          1892 => x"05",
          1893 => x"82",
          1894 => x"90",
          1895 => x"b6",
          1896 => x"05",
          1897 => x"82",
          1898 => x"90",
          1899 => x"b6",
          1900 => x"05",
          1901 => x"ba",
          1902 => x"a4",
          1903 => x"08",
          1904 => x"82",
          1905 => x"f8",
          1906 => x"05",
          1907 => x"08",
          1908 => x"82",
          1909 => x"fc",
          1910 => x"52",
          1911 => x"82",
          1912 => x"fc",
          1913 => x"05",
          1914 => x"08",
          1915 => x"ff",
          1916 => x"b6",
          1917 => x"05",
          1918 => x"b6",
          1919 => x"85",
          1920 => x"b6",
          1921 => x"82",
          1922 => x"02",
          1923 => x"0c",
          1924 => x"82",
          1925 => x"88",
          1926 => x"b6",
          1927 => x"05",
          1928 => x"a4",
          1929 => x"08",
          1930 => x"82",
          1931 => x"fc",
          1932 => x"05",
          1933 => x"08",
          1934 => x"70",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"39",
          1938 => x"08",
          1939 => x"ff",
          1940 => x"a4",
          1941 => x"0c",
          1942 => x"08",
          1943 => x"82",
          1944 => x"88",
          1945 => x"70",
          1946 => x"0c",
          1947 => x"0d",
          1948 => x"0c",
          1949 => x"a4",
          1950 => x"b6",
          1951 => x"3d",
          1952 => x"a4",
          1953 => x"08",
          1954 => x"08",
          1955 => x"82",
          1956 => x"8c",
          1957 => x"71",
          1958 => x"a4",
          1959 => x"08",
          1960 => x"b6",
          1961 => x"05",
          1962 => x"a4",
          1963 => x"08",
          1964 => x"72",
          1965 => x"a4",
          1966 => x"08",
          1967 => x"b6",
          1968 => x"05",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"ff",
          1972 => x"b6",
          1973 => x"05",
          1974 => x"b6",
          1975 => x"84",
          1976 => x"b6",
          1977 => x"82",
          1978 => x"02",
          1979 => x"0c",
          1980 => x"82",
          1981 => x"88",
          1982 => x"b6",
          1983 => x"05",
          1984 => x"a4",
          1985 => x"08",
          1986 => x"08",
          1987 => x"82",
          1988 => x"90",
          1989 => x"2e",
          1990 => x"82",
          1991 => x"90",
          1992 => x"05",
          1993 => x"08",
          1994 => x"82",
          1995 => x"90",
          1996 => x"05",
          1997 => x"08",
          1998 => x"82",
          1999 => x"90",
          2000 => x"2e",
          2001 => x"b6",
          2002 => x"05",
          2003 => x"33",
          2004 => x"08",
          2005 => x"81",
          2006 => x"a4",
          2007 => x"0c",
          2008 => x"08",
          2009 => x"52",
          2010 => x"34",
          2011 => x"08",
          2012 => x"81",
          2013 => x"a4",
          2014 => x"0c",
          2015 => x"82",
          2016 => x"88",
          2017 => x"82",
          2018 => x"51",
          2019 => x"82",
          2020 => x"04",
          2021 => x"08",
          2022 => x"a4",
          2023 => x"0d",
          2024 => x"08",
          2025 => x"80",
          2026 => x"38",
          2027 => x"08",
          2028 => x"52",
          2029 => x"b6",
          2030 => x"05",
          2031 => x"82",
          2032 => x"8c",
          2033 => x"b6",
          2034 => x"05",
          2035 => x"72",
          2036 => x"53",
          2037 => x"71",
          2038 => x"38",
          2039 => x"82",
          2040 => x"88",
          2041 => x"71",
          2042 => x"a4",
          2043 => x"08",
          2044 => x"b6",
          2045 => x"05",
          2046 => x"ff",
          2047 => x"70",
          2048 => x"0b",
          2049 => x"08",
          2050 => x"81",
          2051 => x"b6",
          2052 => x"05",
          2053 => x"82",
          2054 => x"90",
          2055 => x"b6",
          2056 => x"05",
          2057 => x"84",
          2058 => x"39",
          2059 => x"08",
          2060 => x"80",
          2061 => x"38",
          2062 => x"08",
          2063 => x"70",
          2064 => x"70",
          2065 => x"0b",
          2066 => x"08",
          2067 => x"80",
          2068 => x"b6",
          2069 => x"05",
          2070 => x"82",
          2071 => x"8c",
          2072 => x"b6",
          2073 => x"05",
          2074 => x"52",
          2075 => x"38",
          2076 => x"b6",
          2077 => x"05",
          2078 => x"82",
          2079 => x"88",
          2080 => x"33",
          2081 => x"08",
          2082 => x"70",
          2083 => x"31",
          2084 => x"a4",
          2085 => x"0c",
          2086 => x"52",
          2087 => x"80",
          2088 => x"a4",
          2089 => x"0c",
          2090 => x"08",
          2091 => x"82",
          2092 => x"85",
          2093 => x"b6",
          2094 => x"82",
          2095 => x"02",
          2096 => x"0c",
          2097 => x"82",
          2098 => x"88",
          2099 => x"b6",
          2100 => x"05",
          2101 => x"a4",
          2102 => x"08",
          2103 => x"0b",
          2104 => x"08",
          2105 => x"80",
          2106 => x"b6",
          2107 => x"05",
          2108 => x"33",
          2109 => x"08",
          2110 => x"81",
          2111 => x"a4",
          2112 => x"0c",
          2113 => x"06",
          2114 => x"80",
          2115 => x"82",
          2116 => x"8c",
          2117 => x"05",
          2118 => x"08",
          2119 => x"82",
          2120 => x"8c",
          2121 => x"2e",
          2122 => x"be",
          2123 => x"a4",
          2124 => x"08",
          2125 => x"b6",
          2126 => x"05",
          2127 => x"a4",
          2128 => x"08",
          2129 => x"08",
          2130 => x"31",
          2131 => x"a4",
          2132 => x"0c",
          2133 => x"a4",
          2134 => x"08",
          2135 => x"0c",
          2136 => x"82",
          2137 => x"04",
          2138 => x"08",
          2139 => x"a4",
          2140 => x"0d",
          2141 => x"08",
          2142 => x"82",
          2143 => x"fc",
          2144 => x"b6",
          2145 => x"05",
          2146 => x"80",
          2147 => x"b6",
          2148 => x"05",
          2149 => x"82",
          2150 => x"90",
          2151 => x"b6",
          2152 => x"05",
          2153 => x"82",
          2154 => x"90",
          2155 => x"b6",
          2156 => x"05",
          2157 => x"a9",
          2158 => x"a4",
          2159 => x"08",
          2160 => x"b6",
          2161 => x"05",
          2162 => x"71",
          2163 => x"b6",
          2164 => x"05",
          2165 => x"82",
          2166 => x"fc",
          2167 => x"be",
          2168 => x"a4",
          2169 => x"08",
          2170 => x"98",
          2171 => x"3d",
          2172 => x"a4",
          2173 => x"b6",
          2174 => x"82",
          2175 => x"f9",
          2176 => x"0b",
          2177 => x"08",
          2178 => x"82",
          2179 => x"88",
          2180 => x"25",
          2181 => x"b6",
          2182 => x"05",
          2183 => x"b6",
          2184 => x"05",
          2185 => x"82",
          2186 => x"f4",
          2187 => x"b6",
          2188 => x"05",
          2189 => x"81",
          2190 => x"a4",
          2191 => x"0c",
          2192 => x"08",
          2193 => x"82",
          2194 => x"fc",
          2195 => x"b6",
          2196 => x"05",
          2197 => x"b9",
          2198 => x"a4",
          2199 => x"08",
          2200 => x"a4",
          2201 => x"0c",
          2202 => x"b6",
          2203 => x"05",
          2204 => x"a4",
          2205 => x"08",
          2206 => x"0b",
          2207 => x"08",
          2208 => x"82",
          2209 => x"f0",
          2210 => x"b6",
          2211 => x"05",
          2212 => x"82",
          2213 => x"8c",
          2214 => x"82",
          2215 => x"88",
          2216 => x"82",
          2217 => x"b6",
          2218 => x"82",
          2219 => x"f8",
          2220 => x"82",
          2221 => x"fc",
          2222 => x"2e",
          2223 => x"b6",
          2224 => x"05",
          2225 => x"b6",
          2226 => x"05",
          2227 => x"a4",
          2228 => x"08",
          2229 => x"98",
          2230 => x"3d",
          2231 => x"a4",
          2232 => x"b6",
          2233 => x"82",
          2234 => x"fb",
          2235 => x"0b",
          2236 => x"08",
          2237 => x"82",
          2238 => x"88",
          2239 => x"25",
          2240 => x"b6",
          2241 => x"05",
          2242 => x"b6",
          2243 => x"05",
          2244 => x"82",
          2245 => x"fc",
          2246 => x"b6",
          2247 => x"05",
          2248 => x"90",
          2249 => x"a4",
          2250 => x"08",
          2251 => x"a4",
          2252 => x"0c",
          2253 => x"b6",
          2254 => x"05",
          2255 => x"b6",
          2256 => x"05",
          2257 => x"a2",
          2258 => x"98",
          2259 => x"b6",
          2260 => x"05",
          2261 => x"b6",
          2262 => x"05",
          2263 => x"90",
          2264 => x"a4",
          2265 => x"08",
          2266 => x"a4",
          2267 => x"0c",
          2268 => x"08",
          2269 => x"70",
          2270 => x"0c",
          2271 => x"0d",
          2272 => x"0c",
          2273 => x"a4",
          2274 => x"b6",
          2275 => x"3d",
          2276 => x"82",
          2277 => x"8c",
          2278 => x"82",
          2279 => x"88",
          2280 => x"80",
          2281 => x"b6",
          2282 => x"82",
          2283 => x"54",
          2284 => x"82",
          2285 => x"04",
          2286 => x"08",
          2287 => x"a4",
          2288 => x"0d",
          2289 => x"b6",
          2290 => x"05",
          2291 => x"b6",
          2292 => x"05",
          2293 => x"3f",
          2294 => x"08",
          2295 => x"98",
          2296 => x"3d",
          2297 => x"a4",
          2298 => x"b6",
          2299 => x"82",
          2300 => x"fd",
          2301 => x"0b",
          2302 => x"08",
          2303 => x"80",
          2304 => x"a4",
          2305 => x"0c",
          2306 => x"08",
          2307 => x"82",
          2308 => x"88",
          2309 => x"b9",
          2310 => x"a4",
          2311 => x"08",
          2312 => x"38",
          2313 => x"b6",
          2314 => x"05",
          2315 => x"38",
          2316 => x"08",
          2317 => x"10",
          2318 => x"08",
          2319 => x"82",
          2320 => x"fc",
          2321 => x"82",
          2322 => x"fc",
          2323 => x"b8",
          2324 => x"a4",
          2325 => x"08",
          2326 => x"e1",
          2327 => x"a4",
          2328 => x"08",
          2329 => x"08",
          2330 => x"26",
          2331 => x"b6",
          2332 => x"05",
          2333 => x"a4",
          2334 => x"08",
          2335 => x"a4",
          2336 => x"0c",
          2337 => x"08",
          2338 => x"82",
          2339 => x"fc",
          2340 => x"82",
          2341 => x"f8",
          2342 => x"b6",
          2343 => x"05",
          2344 => x"82",
          2345 => x"fc",
          2346 => x"b6",
          2347 => x"05",
          2348 => x"82",
          2349 => x"8c",
          2350 => x"95",
          2351 => x"a4",
          2352 => x"08",
          2353 => x"38",
          2354 => x"08",
          2355 => x"70",
          2356 => x"08",
          2357 => x"51",
          2358 => x"b6",
          2359 => x"05",
          2360 => x"b6",
          2361 => x"05",
          2362 => x"b6",
          2363 => x"05",
          2364 => x"98",
          2365 => x"0d",
          2366 => x"0c",
          2367 => x"a4",
          2368 => x"b6",
          2369 => x"3d",
          2370 => x"82",
          2371 => x"f0",
          2372 => x"b6",
          2373 => x"05",
          2374 => x"73",
          2375 => x"a4",
          2376 => x"08",
          2377 => x"53",
          2378 => x"72",
          2379 => x"08",
          2380 => x"72",
          2381 => x"53",
          2382 => x"09",
          2383 => x"38",
          2384 => x"08",
          2385 => x"70",
          2386 => x"71",
          2387 => x"39",
          2388 => x"08",
          2389 => x"53",
          2390 => x"09",
          2391 => x"38",
          2392 => x"b6",
          2393 => x"05",
          2394 => x"a4",
          2395 => x"08",
          2396 => x"05",
          2397 => x"08",
          2398 => x"33",
          2399 => x"08",
          2400 => x"82",
          2401 => x"f8",
          2402 => x"72",
          2403 => x"81",
          2404 => x"38",
          2405 => x"08",
          2406 => x"70",
          2407 => x"71",
          2408 => x"51",
          2409 => x"82",
          2410 => x"f8",
          2411 => x"b6",
          2412 => x"05",
          2413 => x"a4",
          2414 => x"0c",
          2415 => x"08",
          2416 => x"80",
          2417 => x"38",
          2418 => x"08",
          2419 => x"80",
          2420 => x"38",
          2421 => x"90",
          2422 => x"a4",
          2423 => x"34",
          2424 => x"08",
          2425 => x"70",
          2426 => x"71",
          2427 => x"51",
          2428 => x"82",
          2429 => x"f8",
          2430 => x"a4",
          2431 => x"82",
          2432 => x"f4",
          2433 => x"b6",
          2434 => x"05",
          2435 => x"81",
          2436 => x"70",
          2437 => x"72",
          2438 => x"a4",
          2439 => x"34",
          2440 => x"82",
          2441 => x"f8",
          2442 => x"72",
          2443 => x"38",
          2444 => x"b6",
          2445 => x"05",
          2446 => x"39",
          2447 => x"08",
          2448 => x"53",
          2449 => x"90",
          2450 => x"a4",
          2451 => x"33",
          2452 => x"26",
          2453 => x"39",
          2454 => x"b6",
          2455 => x"05",
          2456 => x"39",
          2457 => x"b6",
          2458 => x"05",
          2459 => x"82",
          2460 => x"f8",
          2461 => x"af",
          2462 => x"38",
          2463 => x"08",
          2464 => x"53",
          2465 => x"83",
          2466 => x"80",
          2467 => x"a4",
          2468 => x"0c",
          2469 => x"8a",
          2470 => x"a4",
          2471 => x"34",
          2472 => x"b6",
          2473 => x"05",
          2474 => x"a4",
          2475 => x"33",
          2476 => x"27",
          2477 => x"82",
          2478 => x"f8",
          2479 => x"80",
          2480 => x"94",
          2481 => x"a4",
          2482 => x"33",
          2483 => x"53",
          2484 => x"a4",
          2485 => x"34",
          2486 => x"08",
          2487 => x"d0",
          2488 => x"72",
          2489 => x"08",
          2490 => x"82",
          2491 => x"f8",
          2492 => x"90",
          2493 => x"38",
          2494 => x"08",
          2495 => x"f9",
          2496 => x"72",
          2497 => x"08",
          2498 => x"82",
          2499 => x"f8",
          2500 => x"72",
          2501 => x"38",
          2502 => x"b6",
          2503 => x"05",
          2504 => x"39",
          2505 => x"08",
          2506 => x"82",
          2507 => x"f4",
          2508 => x"54",
          2509 => x"8d",
          2510 => x"82",
          2511 => x"ec",
          2512 => x"f7",
          2513 => x"a4",
          2514 => x"33",
          2515 => x"a4",
          2516 => x"08",
          2517 => x"a4",
          2518 => x"33",
          2519 => x"b6",
          2520 => x"05",
          2521 => x"a4",
          2522 => x"08",
          2523 => x"05",
          2524 => x"08",
          2525 => x"55",
          2526 => x"82",
          2527 => x"f8",
          2528 => x"a5",
          2529 => x"a4",
          2530 => x"33",
          2531 => x"2e",
          2532 => x"b6",
          2533 => x"05",
          2534 => x"b6",
          2535 => x"05",
          2536 => x"a4",
          2537 => x"08",
          2538 => x"08",
          2539 => x"71",
          2540 => x"0b",
          2541 => x"08",
          2542 => x"82",
          2543 => x"ec",
          2544 => x"b6",
          2545 => x"3d",
          2546 => x"a4",
          2547 => x"b6",
          2548 => x"82",
          2549 => x"f7",
          2550 => x"0b",
          2551 => x"08",
          2552 => x"82",
          2553 => x"8c",
          2554 => x"80",
          2555 => x"b6",
          2556 => x"05",
          2557 => x"51",
          2558 => x"53",
          2559 => x"a4",
          2560 => x"34",
          2561 => x"06",
          2562 => x"2e",
          2563 => x"91",
          2564 => x"a4",
          2565 => x"08",
          2566 => x"05",
          2567 => x"ce",
          2568 => x"a4",
          2569 => x"33",
          2570 => x"2e",
          2571 => x"a4",
          2572 => x"82",
          2573 => x"f0",
          2574 => x"b6",
          2575 => x"05",
          2576 => x"81",
          2577 => x"70",
          2578 => x"72",
          2579 => x"a4",
          2580 => x"34",
          2581 => x"08",
          2582 => x"53",
          2583 => x"09",
          2584 => x"dc",
          2585 => x"a4",
          2586 => x"08",
          2587 => x"05",
          2588 => x"08",
          2589 => x"33",
          2590 => x"08",
          2591 => x"82",
          2592 => x"f8",
          2593 => x"b6",
          2594 => x"05",
          2595 => x"a4",
          2596 => x"08",
          2597 => x"b6",
          2598 => x"a4",
          2599 => x"08",
          2600 => x"84",
          2601 => x"39",
          2602 => x"b6",
          2603 => x"05",
          2604 => x"a4",
          2605 => x"08",
          2606 => x"05",
          2607 => x"08",
          2608 => x"33",
          2609 => x"08",
          2610 => x"81",
          2611 => x"0b",
          2612 => x"08",
          2613 => x"82",
          2614 => x"88",
          2615 => x"08",
          2616 => x"0c",
          2617 => x"53",
          2618 => x"b6",
          2619 => x"05",
          2620 => x"39",
          2621 => x"08",
          2622 => x"53",
          2623 => x"8d",
          2624 => x"82",
          2625 => x"ec",
          2626 => x"80",
          2627 => x"a4",
          2628 => x"33",
          2629 => x"27",
          2630 => x"b6",
          2631 => x"05",
          2632 => x"b9",
          2633 => x"8d",
          2634 => x"82",
          2635 => x"ec",
          2636 => x"d8",
          2637 => x"82",
          2638 => x"f4",
          2639 => x"39",
          2640 => x"08",
          2641 => x"53",
          2642 => x"90",
          2643 => x"a4",
          2644 => x"33",
          2645 => x"26",
          2646 => x"39",
          2647 => x"b6",
          2648 => x"05",
          2649 => x"39",
          2650 => x"b6",
          2651 => x"05",
          2652 => x"82",
          2653 => x"fc",
          2654 => x"b6",
          2655 => x"05",
          2656 => x"73",
          2657 => x"38",
          2658 => x"08",
          2659 => x"53",
          2660 => x"27",
          2661 => x"b6",
          2662 => x"05",
          2663 => x"51",
          2664 => x"b6",
          2665 => x"05",
          2666 => x"a4",
          2667 => x"33",
          2668 => x"53",
          2669 => x"a4",
          2670 => x"34",
          2671 => x"08",
          2672 => x"53",
          2673 => x"ad",
          2674 => x"a4",
          2675 => x"33",
          2676 => x"53",
          2677 => x"a4",
          2678 => x"34",
          2679 => x"08",
          2680 => x"53",
          2681 => x"8d",
          2682 => x"82",
          2683 => x"ec",
          2684 => x"98",
          2685 => x"a4",
          2686 => x"33",
          2687 => x"08",
          2688 => x"54",
          2689 => x"26",
          2690 => x"0b",
          2691 => x"08",
          2692 => x"80",
          2693 => x"b6",
          2694 => x"05",
          2695 => x"b6",
          2696 => x"05",
          2697 => x"b6",
          2698 => x"05",
          2699 => x"82",
          2700 => x"fc",
          2701 => x"b6",
          2702 => x"05",
          2703 => x"81",
          2704 => x"70",
          2705 => x"52",
          2706 => x"33",
          2707 => x"08",
          2708 => x"fe",
          2709 => x"b6",
          2710 => x"05",
          2711 => x"80",
          2712 => x"82",
          2713 => x"fc",
          2714 => x"82",
          2715 => x"fc",
          2716 => x"b6",
          2717 => x"05",
          2718 => x"a4",
          2719 => x"08",
          2720 => x"81",
          2721 => x"a4",
          2722 => x"0c",
          2723 => x"08",
          2724 => x"82",
          2725 => x"8b",
          2726 => x"b6",
          2727 => x"f9",
          2728 => x"70",
          2729 => x"56",
          2730 => x"2e",
          2731 => x"95",
          2732 => x"51",
          2733 => x"82",
          2734 => x"15",
          2735 => x"16",
          2736 => x"cd",
          2737 => x"54",
          2738 => x"09",
          2739 => x"38",
          2740 => x"f1",
          2741 => x"76",
          2742 => x"b1",
          2743 => x"08",
          2744 => x"a3",
          2745 => x"98",
          2746 => x"52",
          2747 => x"e9",
          2748 => x"b6",
          2749 => x"38",
          2750 => x"54",
          2751 => x"ff",
          2752 => x"17",
          2753 => x"06",
          2754 => x"77",
          2755 => x"ff",
          2756 => x"b6",
          2757 => x"3d",
          2758 => x"3d",
          2759 => x"71",
          2760 => x"8e",
          2761 => x"29",
          2762 => x"05",
          2763 => x"04",
          2764 => x"51",
          2765 => x"82",
          2766 => x"80",
          2767 => x"9b",
          2768 => x"f2",
          2769 => x"c4",
          2770 => x"39",
          2771 => x"51",
          2772 => x"82",
          2773 => x"80",
          2774 => x"9b",
          2775 => x"d6",
          2776 => x"88",
          2777 => x"39",
          2778 => x"51",
          2779 => x"82",
          2780 => x"80",
          2781 => x"9c",
          2782 => x"39",
          2783 => x"51",
          2784 => x"9d",
          2785 => x"39",
          2786 => x"51",
          2787 => x"9d",
          2788 => x"39",
          2789 => x"51",
          2790 => x"9d",
          2791 => x"39",
          2792 => x"51",
          2793 => x"9e",
          2794 => x"39",
          2795 => x"51",
          2796 => x"9e",
          2797 => x"ad",
          2798 => x"0d",
          2799 => x"0d",
          2800 => x"56",
          2801 => x"26",
          2802 => x"52",
          2803 => x"29",
          2804 => x"87",
          2805 => x"51",
          2806 => x"82",
          2807 => x"52",
          2808 => x"a1",
          2809 => x"98",
          2810 => x"53",
          2811 => x"9e",
          2812 => x"bb",
          2813 => x"3d",
          2814 => x"3d",
          2815 => x"84",
          2816 => x"05",
          2817 => x"80",
          2818 => x"70",
          2819 => x"25",
          2820 => x"59",
          2821 => x"87",
          2822 => x"38",
          2823 => x"76",
          2824 => x"ff",
          2825 => x"93",
          2826 => x"82",
          2827 => x"76",
          2828 => x"70",
          2829 => x"ff",
          2830 => x"b6",
          2831 => x"82",
          2832 => x"b9",
          2833 => x"98",
          2834 => x"98",
          2835 => x"b6",
          2836 => x"96",
          2837 => x"54",
          2838 => x"77",
          2839 => x"81",
          2840 => x"82",
          2841 => x"57",
          2842 => x"08",
          2843 => x"55",
          2844 => x"89",
          2845 => x"75",
          2846 => x"d7",
          2847 => x"d8",
          2848 => x"8c",
          2849 => x"30",
          2850 => x"80",
          2851 => x"70",
          2852 => x"06",
          2853 => x"56",
          2854 => x"90",
          2855 => x"f0",
          2856 => x"98",
          2857 => x"78",
          2858 => x"3f",
          2859 => x"82",
          2860 => x"96",
          2861 => x"f7",
          2862 => x"02",
          2863 => x"05",
          2864 => x"ff",
          2865 => x"7c",
          2866 => x"fe",
          2867 => x"b6",
          2868 => x"cb",
          2869 => x"2e",
          2870 => x"81",
          2871 => x"bf",
          2872 => x"e8",
          2873 => x"e8",
          2874 => x"e8",
          2875 => x"f0",
          2876 => x"cd",
          2877 => x"82",
          2878 => x"52",
          2879 => x"51",
          2880 => x"3f",
          2881 => x"56",
          2882 => x"54",
          2883 => x"53",
          2884 => x"51",
          2885 => x"b6",
          2886 => x"83",
          2887 => x"78",
          2888 => x"0c",
          2889 => x"04",
          2890 => x"7f",
          2891 => x"8c",
          2892 => x"05",
          2893 => x"15",
          2894 => x"5c",
          2895 => x"5e",
          2896 => x"9f",
          2897 => x"b9",
          2898 => x"9f",
          2899 => x"b9",
          2900 => x"55",
          2901 => x"81",
          2902 => x"90",
          2903 => x"7b",
          2904 => x"38",
          2905 => x"74",
          2906 => x"7a",
          2907 => x"72",
          2908 => x"9f",
          2909 => x"b8",
          2910 => x"39",
          2911 => x"51",
          2912 => x"3f",
          2913 => x"80",
          2914 => x"18",
          2915 => x"27",
          2916 => x"08",
          2917 => x"ac",
          2918 => x"be",
          2919 => x"82",
          2920 => x"ff",
          2921 => x"84",
          2922 => x"39",
          2923 => x"72",
          2924 => x"38",
          2925 => x"82",
          2926 => x"ff",
          2927 => x"89",
          2928 => x"d4",
          2929 => x"92",
          2930 => x"55",
          2931 => x"08",
          2932 => x"d7",
          2933 => x"fc",
          2934 => x"d8",
          2935 => x"fa",
          2936 => x"74",
          2937 => x"c6",
          2938 => x"70",
          2939 => x"80",
          2940 => x"27",
          2941 => x"56",
          2942 => x"74",
          2943 => x"81",
          2944 => x"06",
          2945 => x"06",
          2946 => x"80",
          2947 => x"73",
          2948 => x"8a",
          2949 => x"ec",
          2950 => x"51",
          2951 => x"cd",
          2952 => x"a0",
          2953 => x"3f",
          2954 => x"ff",
          2955 => x"9f",
          2956 => x"b1",
          2957 => x"79",
          2958 => x"9c",
          2959 => x"b6",
          2960 => x"2b",
          2961 => x"51",
          2962 => x"2e",
          2963 => x"aa",
          2964 => x"3f",
          2965 => x"08",
          2966 => x"98",
          2967 => x"32",
          2968 => x"9b",
          2969 => x"70",
          2970 => x"75",
          2971 => x"58",
          2972 => x"51",
          2973 => x"24",
          2974 => x"9b",
          2975 => x"06",
          2976 => x"53",
          2977 => x"1e",
          2978 => x"26",
          2979 => x"ff",
          2980 => x"b6",
          2981 => x"3d",
          2982 => x"3d",
          2983 => x"05",
          2984 => x"e0",
          2985 => x"e4",
          2986 => x"b6",
          2987 => x"b4",
          2988 => x"a5",
          2989 => x"9f",
          2990 => x"9f",
          2991 => x"b4",
          2992 => x"82",
          2993 => x"ff",
          2994 => x"74",
          2995 => x"38",
          2996 => x"86",
          2997 => x"fe",
          2998 => x"c0",
          2999 => x"53",
          3000 => x"81",
          3001 => x"3f",
          3002 => x"51",
          3003 => x"80",
          3004 => x"3f",
          3005 => x"70",
          3006 => x"52",
          3007 => x"92",
          3008 => x"97",
          3009 => x"a0",
          3010 => x"85",
          3011 => x"97",
          3012 => x"82",
          3013 => x"06",
          3014 => x"80",
          3015 => x"81",
          3016 => x"3f",
          3017 => x"51",
          3018 => x"80",
          3019 => x"3f",
          3020 => x"70",
          3021 => x"52",
          3022 => x"92",
          3023 => x"97",
          3024 => x"a0",
          3025 => x"c9",
          3026 => x"97",
          3027 => x"84",
          3028 => x"06",
          3029 => x"80",
          3030 => x"81",
          3031 => x"3f",
          3032 => x"51",
          3033 => x"80",
          3034 => x"3f",
          3035 => x"70",
          3036 => x"52",
          3037 => x"92",
          3038 => x"96",
          3039 => x"a1",
          3040 => x"8d",
          3041 => x"96",
          3042 => x"86",
          3043 => x"06",
          3044 => x"80",
          3045 => x"81",
          3046 => x"3f",
          3047 => x"51",
          3048 => x"80",
          3049 => x"3f",
          3050 => x"70",
          3051 => x"52",
          3052 => x"92",
          3053 => x"96",
          3054 => x"a1",
          3055 => x"d1",
          3056 => x"96",
          3057 => x"88",
          3058 => x"06",
          3059 => x"80",
          3060 => x"81",
          3061 => x"3f",
          3062 => x"51",
          3063 => x"80",
          3064 => x"3f",
          3065 => x"84",
          3066 => x"fb",
          3067 => x"02",
          3068 => x"05",
          3069 => x"56",
          3070 => x"75",
          3071 => x"3f",
          3072 => x"b1",
          3073 => x"73",
          3074 => x"53",
          3075 => x"52",
          3076 => x"51",
          3077 => x"3f",
          3078 => x"08",
          3079 => x"b6",
          3080 => x"80",
          3081 => x"31",
          3082 => x"73",
          3083 => x"b1",
          3084 => x"0b",
          3085 => x"33",
          3086 => x"2e",
          3087 => x"af",
          3088 => x"98",
          3089 => x"75",
          3090 => x"ba",
          3091 => x"98",
          3092 => x"8b",
          3093 => x"98",
          3094 => x"89",
          3095 => x"82",
          3096 => x"81",
          3097 => x"82",
          3098 => x"82",
          3099 => x"0b",
          3100 => x"94",
          3101 => x"82",
          3102 => x"06",
          3103 => x"a2",
          3104 => x"52",
          3105 => x"bc",
          3106 => x"82",
          3107 => x"87",
          3108 => x"ce",
          3109 => x"70",
          3110 => x"94",
          3111 => x"81",
          3112 => x"80",
          3113 => x"82",
          3114 => x"81",
          3115 => x"78",
          3116 => x"81",
          3117 => x"96",
          3118 => x"53",
          3119 => x"52",
          3120 => x"a3",
          3121 => x"78",
          3122 => x"c4",
          3123 => x"ef",
          3124 => x"98",
          3125 => x"88",
          3126 => x"94",
          3127 => x"39",
          3128 => x"5d",
          3129 => x"51",
          3130 => x"3f",
          3131 => x"46",
          3132 => x"52",
          3133 => x"f3",
          3134 => x"ff",
          3135 => x"f3",
          3136 => x"b6",
          3137 => x"2b",
          3138 => x"51",
          3139 => x"c2",
          3140 => x"38",
          3141 => x"24",
          3142 => x"bd",
          3143 => x"38",
          3144 => x"90",
          3145 => x"2e",
          3146 => x"78",
          3147 => x"da",
          3148 => x"39",
          3149 => x"2e",
          3150 => x"78",
          3151 => x"85",
          3152 => x"bf",
          3153 => x"38",
          3154 => x"78",
          3155 => x"89",
          3156 => x"80",
          3157 => x"38",
          3158 => x"2e",
          3159 => x"78",
          3160 => x"89",
          3161 => x"9f",
          3162 => x"83",
          3163 => x"38",
          3164 => x"24",
          3165 => x"81",
          3166 => x"eb",
          3167 => x"39",
          3168 => x"2e",
          3169 => x"89",
          3170 => x"3d",
          3171 => x"53",
          3172 => x"51",
          3173 => x"82",
          3174 => x"80",
          3175 => x"38",
          3176 => x"fc",
          3177 => x"84",
          3178 => x"a2",
          3179 => x"98",
          3180 => x"fe",
          3181 => x"3d",
          3182 => x"53",
          3183 => x"51",
          3184 => x"82",
          3185 => x"86",
          3186 => x"98",
          3187 => x"a2",
          3188 => x"b0",
          3189 => x"63",
          3190 => x"7b",
          3191 => x"38",
          3192 => x"7a",
          3193 => x"5c",
          3194 => x"26",
          3195 => x"db",
          3196 => x"ff",
          3197 => x"ff",
          3198 => x"eb",
          3199 => x"b6",
          3200 => x"2e",
          3201 => x"b4",
          3202 => x"11",
          3203 => x"05",
          3204 => x"3f",
          3205 => x"08",
          3206 => x"c8",
          3207 => x"fe",
          3208 => x"ff",
          3209 => x"eb",
          3210 => x"b6",
          3211 => x"2e",
          3212 => x"82",
          3213 => x"ff",
          3214 => x"63",
          3215 => x"27",
          3216 => x"61",
          3217 => x"81",
          3218 => x"79",
          3219 => x"05",
          3220 => x"b4",
          3221 => x"11",
          3222 => x"05",
          3223 => x"3f",
          3224 => x"08",
          3225 => x"fc",
          3226 => x"fe",
          3227 => x"ff",
          3228 => x"ea",
          3229 => x"b6",
          3230 => x"2e",
          3231 => x"b4",
          3232 => x"11",
          3233 => x"05",
          3234 => x"3f",
          3235 => x"08",
          3236 => x"d0",
          3237 => x"ec",
          3238 => x"be",
          3239 => x"79",
          3240 => x"38",
          3241 => x"7b",
          3242 => x"5b",
          3243 => x"92",
          3244 => x"7a",
          3245 => x"53",
          3246 => x"a2",
          3247 => x"ae",
          3248 => x"1a",
          3249 => x"43",
          3250 => x"8a",
          3251 => x"3f",
          3252 => x"b4",
          3253 => x"11",
          3254 => x"05",
          3255 => x"3f",
          3256 => x"08",
          3257 => x"82",
          3258 => x"59",
          3259 => x"89",
          3260 => x"bc",
          3261 => x"cd",
          3262 => x"85",
          3263 => x"80",
          3264 => x"82",
          3265 => x"44",
          3266 => x"b5",
          3267 => x"78",
          3268 => x"38",
          3269 => x"08",
          3270 => x"82",
          3271 => x"59",
          3272 => x"88",
          3273 => x"d4",
          3274 => x"39",
          3275 => x"33",
          3276 => x"2e",
          3277 => x"b4",
          3278 => x"89",
          3279 => x"ec",
          3280 => x"05",
          3281 => x"fe",
          3282 => x"ff",
          3283 => x"e8",
          3284 => x"b6",
          3285 => x"de",
          3286 => x"84",
          3287 => x"80",
          3288 => x"82",
          3289 => x"43",
          3290 => x"82",
          3291 => x"59",
          3292 => x"88",
          3293 => x"c8",
          3294 => x"39",
          3295 => x"33",
          3296 => x"2e",
          3297 => x"b4",
          3298 => x"aa",
          3299 => x"87",
          3300 => x"80",
          3301 => x"82",
          3302 => x"43",
          3303 => x"b5",
          3304 => x"78",
          3305 => x"38",
          3306 => x"08",
          3307 => x"82",
          3308 => x"88",
          3309 => x"3d",
          3310 => x"53",
          3311 => x"51",
          3312 => x"82",
          3313 => x"80",
          3314 => x"80",
          3315 => x"7a",
          3316 => x"38",
          3317 => x"90",
          3318 => x"70",
          3319 => x"2a",
          3320 => x"51",
          3321 => x"78",
          3322 => x"38",
          3323 => x"83",
          3324 => x"82",
          3325 => x"c7",
          3326 => x"55",
          3327 => x"53",
          3328 => x"51",
          3329 => x"82",
          3330 => x"86",
          3331 => x"3d",
          3332 => x"53",
          3333 => x"51",
          3334 => x"82",
          3335 => x"80",
          3336 => x"38",
          3337 => x"fc",
          3338 => x"84",
          3339 => x"9e",
          3340 => x"98",
          3341 => x"a4",
          3342 => x"02",
          3343 => x"33",
          3344 => x"81",
          3345 => x"3d",
          3346 => x"53",
          3347 => x"51",
          3348 => x"82",
          3349 => x"e1",
          3350 => x"39",
          3351 => x"54",
          3352 => x"b0",
          3353 => x"f2",
          3354 => x"e8",
          3355 => x"f8",
          3356 => x"ff",
          3357 => x"79",
          3358 => x"59",
          3359 => x"f8",
          3360 => x"79",
          3361 => x"b4",
          3362 => x"11",
          3363 => x"05",
          3364 => x"3f",
          3365 => x"08",
          3366 => x"38",
          3367 => x"80",
          3368 => x"79",
          3369 => x"05",
          3370 => x"39",
          3371 => x"51",
          3372 => x"ff",
          3373 => x"3d",
          3374 => x"53",
          3375 => x"51",
          3376 => x"82",
          3377 => x"80",
          3378 => x"38",
          3379 => x"f0",
          3380 => x"84",
          3381 => x"a5",
          3382 => x"98",
          3383 => x"a5",
          3384 => x"02",
          3385 => x"79",
          3386 => x"5b",
          3387 => x"b4",
          3388 => x"11",
          3389 => x"05",
          3390 => x"3f",
          3391 => x"08",
          3392 => x"e0",
          3393 => x"22",
          3394 => x"a3",
          3395 => x"a9",
          3396 => x"cd",
          3397 => x"80",
          3398 => x"51",
          3399 => x"3f",
          3400 => x"33",
          3401 => x"2e",
          3402 => x"78",
          3403 => x"38",
          3404 => x"41",
          3405 => x"3d",
          3406 => x"53",
          3407 => x"51",
          3408 => x"82",
          3409 => x"80",
          3410 => x"60",
          3411 => x"05",
          3412 => x"82",
          3413 => x"78",
          3414 => x"39",
          3415 => x"51",
          3416 => x"ff",
          3417 => x"3d",
          3418 => x"53",
          3419 => x"51",
          3420 => x"82",
          3421 => x"80",
          3422 => x"38",
          3423 => x"f0",
          3424 => x"84",
          3425 => x"f5",
          3426 => x"98",
          3427 => x"a0",
          3428 => x"71",
          3429 => x"84",
          3430 => x"3d",
          3431 => x"53",
          3432 => x"51",
          3433 => x"82",
          3434 => x"e5",
          3435 => x"39",
          3436 => x"54",
          3437 => x"cc",
          3438 => x"9e",
          3439 => x"e8",
          3440 => x"f8",
          3441 => x"ff",
          3442 => x"79",
          3443 => x"59",
          3444 => x"f6",
          3445 => x"79",
          3446 => x"b4",
          3447 => x"11",
          3448 => x"05",
          3449 => x"3f",
          3450 => x"08",
          3451 => x"38",
          3452 => x"0c",
          3453 => x"05",
          3454 => x"39",
          3455 => x"51",
          3456 => x"ff",
          3457 => x"3d",
          3458 => x"53",
          3459 => x"51",
          3460 => x"82",
          3461 => x"80",
          3462 => x"38",
          3463 => x"a3",
          3464 => x"a7",
          3465 => x"59",
          3466 => x"3d",
          3467 => x"53",
          3468 => x"51",
          3469 => x"82",
          3470 => x"80",
          3471 => x"38",
          3472 => x"a3",
          3473 => x"a7",
          3474 => x"59",
          3475 => x"b6",
          3476 => x"2e",
          3477 => x"82",
          3478 => x"52",
          3479 => x"51",
          3480 => x"3f",
          3481 => x"82",
          3482 => x"c2",
          3483 => x"a6",
          3484 => x"f0",
          3485 => x"cc",
          3486 => x"3f",
          3487 => x"a8",
          3488 => x"3f",
          3489 => x"79",
          3490 => x"59",
          3491 => x"f4",
          3492 => x"7d",
          3493 => x"80",
          3494 => x"38",
          3495 => x"84",
          3496 => x"ca",
          3497 => x"98",
          3498 => x"5b",
          3499 => x"b2",
          3500 => x"24",
          3501 => x"81",
          3502 => x"80",
          3503 => x"83",
          3504 => x"80",
          3505 => x"a4",
          3506 => x"55",
          3507 => x"54",
          3508 => x"a4",
          3509 => x"3d",
          3510 => x"51",
          3511 => x"3f",
          3512 => x"52",
          3513 => x"b0",
          3514 => x"89",
          3515 => x"7b",
          3516 => x"e4",
          3517 => x"82",
          3518 => x"b4",
          3519 => x"05",
          3520 => x"be",
          3521 => x"7b",
          3522 => x"82",
          3523 => x"b4",
          3524 => x"05",
          3525 => x"aa",
          3526 => x"bc",
          3527 => x"c8",
          3528 => x"64",
          3529 => x"82",
          3530 => x"82",
          3531 => x"b4",
          3532 => x"05",
          3533 => x"3f",
          3534 => x"08",
          3535 => x"08",
          3536 => x"70",
          3537 => x"25",
          3538 => x"5f",
          3539 => x"83",
          3540 => x"81",
          3541 => x"06",
          3542 => x"2e",
          3543 => x"1b",
          3544 => x"06",
          3545 => x"fe",
          3546 => x"81",
          3547 => x"32",
          3548 => x"8a",
          3549 => x"2e",
          3550 => x"f2",
          3551 => x"a5",
          3552 => x"e1",
          3553 => x"39",
          3554 => x"80",
          3555 => x"c8",
          3556 => x"94",
          3557 => x"54",
          3558 => x"80",
          3559 => x"d7",
          3560 => x"b6",
          3561 => x"2b",
          3562 => x"53",
          3563 => x"52",
          3564 => x"d1",
          3565 => x"b6",
          3566 => x"75",
          3567 => x"94",
          3568 => x"54",
          3569 => x"80",
          3570 => x"d7",
          3571 => x"b6",
          3572 => x"2b",
          3573 => x"53",
          3574 => x"52",
          3575 => x"a5",
          3576 => x"b6",
          3577 => x"75",
          3578 => x"83",
          3579 => x"94",
          3580 => x"80",
          3581 => x"c0",
          3582 => x"80",
          3583 => x"80",
          3584 => x"83",
          3585 => x"99",
          3586 => x"5c",
          3587 => x"0b",
          3588 => x"88",
          3589 => x"72",
          3590 => x"ec",
          3591 => x"be",
          3592 => x"3f",
          3593 => x"51",
          3594 => x"3f",
          3595 => x"51",
          3596 => x"3f",
          3597 => x"51",
          3598 => x"81",
          3599 => x"3f",
          3600 => x"80",
          3601 => x"0d",
          3602 => x"53",
          3603 => x"52",
          3604 => x"82",
          3605 => x"81",
          3606 => x"07",
          3607 => x"52",
          3608 => x"e8",
          3609 => x"b6",
          3610 => x"3d",
          3611 => x"3d",
          3612 => x"08",
          3613 => x"73",
          3614 => x"74",
          3615 => x"38",
          3616 => x"70",
          3617 => x"81",
          3618 => x"81",
          3619 => x"39",
          3620 => x"70",
          3621 => x"81",
          3622 => x"81",
          3623 => x"54",
          3624 => x"81",
          3625 => x"06",
          3626 => x"39",
          3627 => x"80",
          3628 => x"54",
          3629 => x"83",
          3630 => x"70",
          3631 => x"38",
          3632 => x"98",
          3633 => x"52",
          3634 => x"52",
          3635 => x"2e",
          3636 => x"54",
          3637 => x"84",
          3638 => x"38",
          3639 => x"52",
          3640 => x"2e",
          3641 => x"83",
          3642 => x"70",
          3643 => x"30",
          3644 => x"76",
          3645 => x"51",
          3646 => x"88",
          3647 => x"70",
          3648 => x"34",
          3649 => x"72",
          3650 => x"b6",
          3651 => x"3d",
          3652 => x"3d",
          3653 => x"72",
          3654 => x"91",
          3655 => x"fc",
          3656 => x"51",
          3657 => x"82",
          3658 => x"85",
          3659 => x"83",
          3660 => x"72",
          3661 => x"0c",
          3662 => x"04",
          3663 => x"76",
          3664 => x"ff",
          3665 => x"81",
          3666 => x"26",
          3667 => x"83",
          3668 => x"05",
          3669 => x"70",
          3670 => x"8a",
          3671 => x"33",
          3672 => x"70",
          3673 => x"fe",
          3674 => x"33",
          3675 => x"70",
          3676 => x"f2",
          3677 => x"33",
          3678 => x"70",
          3679 => x"e6",
          3680 => x"22",
          3681 => x"74",
          3682 => x"80",
          3683 => x"13",
          3684 => x"52",
          3685 => x"26",
          3686 => x"81",
          3687 => x"98",
          3688 => x"22",
          3689 => x"bc",
          3690 => x"33",
          3691 => x"b8",
          3692 => x"33",
          3693 => x"b4",
          3694 => x"33",
          3695 => x"b0",
          3696 => x"33",
          3697 => x"ac",
          3698 => x"33",
          3699 => x"a8",
          3700 => x"c0",
          3701 => x"73",
          3702 => x"a0",
          3703 => x"87",
          3704 => x"0c",
          3705 => x"82",
          3706 => x"86",
          3707 => x"f3",
          3708 => x"5b",
          3709 => x"9c",
          3710 => x"0c",
          3711 => x"bc",
          3712 => x"7b",
          3713 => x"98",
          3714 => x"79",
          3715 => x"87",
          3716 => x"08",
          3717 => x"1c",
          3718 => x"98",
          3719 => x"79",
          3720 => x"87",
          3721 => x"08",
          3722 => x"1c",
          3723 => x"98",
          3724 => x"79",
          3725 => x"87",
          3726 => x"08",
          3727 => x"1c",
          3728 => x"98",
          3729 => x"79",
          3730 => x"80",
          3731 => x"83",
          3732 => x"59",
          3733 => x"ff",
          3734 => x"1b",
          3735 => x"1b",
          3736 => x"1b",
          3737 => x"1b",
          3738 => x"1b",
          3739 => x"83",
          3740 => x"52",
          3741 => x"51",
          3742 => x"3f",
          3743 => x"04",
          3744 => x"02",
          3745 => x"82",
          3746 => x"70",
          3747 => x"58",
          3748 => x"c0",
          3749 => x"75",
          3750 => x"38",
          3751 => x"94",
          3752 => x"70",
          3753 => x"81",
          3754 => x"52",
          3755 => x"8c",
          3756 => x"2a",
          3757 => x"51",
          3758 => x"38",
          3759 => x"70",
          3760 => x"51",
          3761 => x"8d",
          3762 => x"2a",
          3763 => x"51",
          3764 => x"be",
          3765 => x"ff",
          3766 => x"c0",
          3767 => x"70",
          3768 => x"38",
          3769 => x"90",
          3770 => x"0c",
          3771 => x"98",
          3772 => x"0d",
          3773 => x"0d",
          3774 => x"33",
          3775 => x"9f",
          3776 => x"52",
          3777 => x"b8",
          3778 => x"0d",
          3779 => x"0d",
          3780 => x"33",
          3781 => x"2e",
          3782 => x"87",
          3783 => x"8d",
          3784 => x"82",
          3785 => x"70",
          3786 => x"58",
          3787 => x"94",
          3788 => x"80",
          3789 => x"87",
          3790 => x"53",
          3791 => x"96",
          3792 => x"06",
          3793 => x"72",
          3794 => x"38",
          3795 => x"70",
          3796 => x"53",
          3797 => x"74",
          3798 => x"81",
          3799 => x"72",
          3800 => x"38",
          3801 => x"70",
          3802 => x"53",
          3803 => x"38",
          3804 => x"06",
          3805 => x"94",
          3806 => x"80",
          3807 => x"87",
          3808 => x"54",
          3809 => x"80",
          3810 => x"98",
          3811 => x"0d",
          3812 => x"0d",
          3813 => x"74",
          3814 => x"ff",
          3815 => x"57",
          3816 => x"80",
          3817 => x"81",
          3818 => x"15",
          3819 => x"33",
          3820 => x"06",
          3821 => x"58",
          3822 => x"84",
          3823 => x"2e",
          3824 => x"c0",
          3825 => x"70",
          3826 => x"2a",
          3827 => x"53",
          3828 => x"80",
          3829 => x"71",
          3830 => x"81",
          3831 => x"70",
          3832 => x"81",
          3833 => x"06",
          3834 => x"80",
          3835 => x"71",
          3836 => x"81",
          3837 => x"70",
          3838 => x"74",
          3839 => x"51",
          3840 => x"80",
          3841 => x"2e",
          3842 => x"c0",
          3843 => x"77",
          3844 => x"17",
          3845 => x"81",
          3846 => x"53",
          3847 => x"86",
          3848 => x"b6",
          3849 => x"3d",
          3850 => x"3d",
          3851 => x"b8",
          3852 => x"ff",
          3853 => x"87",
          3854 => x"51",
          3855 => x"86",
          3856 => x"94",
          3857 => x"08",
          3858 => x"70",
          3859 => x"51",
          3860 => x"2e",
          3861 => x"81",
          3862 => x"87",
          3863 => x"52",
          3864 => x"86",
          3865 => x"94",
          3866 => x"08",
          3867 => x"06",
          3868 => x"0c",
          3869 => x"0d",
          3870 => x"3f",
          3871 => x"08",
          3872 => x"82",
          3873 => x"04",
          3874 => x"82",
          3875 => x"70",
          3876 => x"52",
          3877 => x"94",
          3878 => x"80",
          3879 => x"87",
          3880 => x"52",
          3881 => x"82",
          3882 => x"06",
          3883 => x"ff",
          3884 => x"2e",
          3885 => x"81",
          3886 => x"87",
          3887 => x"52",
          3888 => x"86",
          3889 => x"94",
          3890 => x"08",
          3891 => x"70",
          3892 => x"53",
          3893 => x"b6",
          3894 => x"3d",
          3895 => x"3d",
          3896 => x"9e",
          3897 => x"9c",
          3898 => x"51",
          3899 => x"2e",
          3900 => x"87",
          3901 => x"08",
          3902 => x"0c",
          3903 => x"a8",
          3904 => x"c0",
          3905 => x"9e",
          3906 => x"b4",
          3907 => x"c0",
          3908 => x"82",
          3909 => x"87",
          3910 => x"08",
          3911 => x"0c",
          3912 => x"a0",
          3913 => x"d0",
          3914 => x"9e",
          3915 => x"b4",
          3916 => x"c0",
          3917 => x"82",
          3918 => x"87",
          3919 => x"08",
          3920 => x"0c",
          3921 => x"b8",
          3922 => x"e0",
          3923 => x"9e",
          3924 => x"b4",
          3925 => x"c0",
          3926 => x"82",
          3927 => x"87",
          3928 => x"08",
          3929 => x"0c",
          3930 => x"80",
          3931 => x"82",
          3932 => x"87",
          3933 => x"08",
          3934 => x"0c",
          3935 => x"88",
          3936 => x"f8",
          3937 => x"9e",
          3938 => x"b4",
          3939 => x"0b",
          3940 => x"34",
          3941 => x"c0",
          3942 => x"70",
          3943 => x"06",
          3944 => x"70",
          3945 => x"38",
          3946 => x"82",
          3947 => x"80",
          3948 => x"9e",
          3949 => x"88",
          3950 => x"51",
          3951 => x"80",
          3952 => x"81",
          3953 => x"b5",
          3954 => x"0b",
          3955 => x"90",
          3956 => x"80",
          3957 => x"52",
          3958 => x"2e",
          3959 => x"52",
          3960 => x"83",
          3961 => x"87",
          3962 => x"08",
          3963 => x"80",
          3964 => x"52",
          3965 => x"83",
          3966 => x"71",
          3967 => x"34",
          3968 => x"c0",
          3969 => x"70",
          3970 => x"06",
          3971 => x"70",
          3972 => x"38",
          3973 => x"82",
          3974 => x"80",
          3975 => x"9e",
          3976 => x"90",
          3977 => x"51",
          3978 => x"80",
          3979 => x"81",
          3980 => x"b5",
          3981 => x"0b",
          3982 => x"90",
          3983 => x"80",
          3984 => x"52",
          3985 => x"2e",
          3986 => x"52",
          3987 => x"87",
          3988 => x"87",
          3989 => x"08",
          3990 => x"80",
          3991 => x"52",
          3992 => x"83",
          3993 => x"71",
          3994 => x"34",
          3995 => x"c0",
          3996 => x"70",
          3997 => x"06",
          3998 => x"70",
          3999 => x"38",
          4000 => x"82",
          4001 => x"80",
          4002 => x"9e",
          4003 => x"80",
          4004 => x"51",
          4005 => x"80",
          4006 => x"81",
          4007 => x"b5",
          4008 => x"0b",
          4009 => x"90",
          4010 => x"80",
          4011 => x"52",
          4012 => x"83",
          4013 => x"71",
          4014 => x"34",
          4015 => x"90",
          4016 => x"80",
          4017 => x"2a",
          4018 => x"70",
          4019 => x"34",
          4020 => x"c0",
          4021 => x"70",
          4022 => x"51",
          4023 => x"80",
          4024 => x"81",
          4025 => x"b5",
          4026 => x"c0",
          4027 => x"70",
          4028 => x"70",
          4029 => x"51",
          4030 => x"b5",
          4031 => x"0b",
          4032 => x"90",
          4033 => x"06",
          4034 => x"70",
          4035 => x"38",
          4036 => x"82",
          4037 => x"87",
          4038 => x"08",
          4039 => x"51",
          4040 => x"b5",
          4041 => x"3d",
          4042 => x"3d",
          4043 => x"d8",
          4044 => x"a6",
          4045 => x"80",
          4046 => x"80",
          4047 => x"82",
          4048 => x"ff",
          4049 => x"82",
          4050 => x"ff",
          4051 => x"82",
          4052 => x"54",
          4053 => x"94",
          4054 => x"dc",
          4055 => x"e0",
          4056 => x"52",
          4057 => x"51",
          4058 => x"3f",
          4059 => x"33",
          4060 => x"2e",
          4061 => x"b4",
          4062 => x"b4",
          4063 => x"54",
          4064 => x"b4",
          4065 => x"d2",
          4066 => x"84",
          4067 => x"80",
          4068 => x"82",
          4069 => x"82",
          4070 => x"11",
          4071 => x"a6",
          4072 => x"94",
          4073 => x"b5",
          4074 => x"73",
          4075 => x"38",
          4076 => x"08",
          4077 => x"08",
          4078 => x"82",
          4079 => x"ff",
          4080 => x"82",
          4081 => x"54",
          4082 => x"94",
          4083 => x"cc",
          4084 => x"d0",
          4085 => x"52",
          4086 => x"51",
          4087 => x"3f",
          4088 => x"33",
          4089 => x"2e",
          4090 => x"b5",
          4091 => x"82",
          4092 => x"ff",
          4093 => x"82",
          4094 => x"54",
          4095 => x"8e",
          4096 => x"90",
          4097 => x"a7",
          4098 => x"93",
          4099 => x"b5",
          4100 => x"73",
          4101 => x"38",
          4102 => x"33",
          4103 => x"e4",
          4104 => x"b6",
          4105 => x"81",
          4106 => x"80",
          4107 => x"82",
          4108 => x"ff",
          4109 => x"82",
          4110 => x"54",
          4111 => x"89",
          4112 => x"98",
          4113 => x"9d",
          4114 => x"88",
          4115 => x"80",
          4116 => x"82",
          4117 => x"ff",
          4118 => x"82",
          4119 => x"54",
          4120 => x"89",
          4121 => x"b0",
          4122 => x"f9",
          4123 => x"8a",
          4124 => x"80",
          4125 => x"82",
          4126 => x"ff",
          4127 => x"82",
          4128 => x"ff",
          4129 => x"82",
          4130 => x"52",
          4131 => x"51",
          4132 => x"3f",
          4133 => x"08",
          4134 => x"f4",
          4135 => x"ba",
          4136 => x"ec",
          4137 => x"a9",
          4138 => x"92",
          4139 => x"a9",
          4140 => x"ae",
          4141 => x"b4",
          4142 => x"82",
          4143 => x"ff",
          4144 => x"82",
          4145 => x"56",
          4146 => x"52",
          4147 => x"b5",
          4148 => x"98",
          4149 => x"c0",
          4150 => x"31",
          4151 => x"b6",
          4152 => x"82",
          4153 => x"ff",
          4154 => x"82",
          4155 => x"54",
          4156 => x"a9",
          4157 => x"f8",
          4158 => x"84",
          4159 => x"51",
          4160 => x"82",
          4161 => x"bd",
          4162 => x"76",
          4163 => x"54",
          4164 => x"08",
          4165 => x"a0",
          4166 => x"be",
          4167 => x"82",
          4168 => x"80",
          4169 => x"82",
          4170 => x"56",
          4171 => x"52",
          4172 => x"d1",
          4173 => x"98",
          4174 => x"c0",
          4175 => x"31",
          4176 => x"b6",
          4177 => x"82",
          4178 => x"ff",
          4179 => x"8a",
          4180 => x"b3",
          4181 => x"0d",
          4182 => x"0d",
          4183 => x"33",
          4184 => x"71",
          4185 => x"38",
          4186 => x"82",
          4187 => x"52",
          4188 => x"82",
          4189 => x"9d",
          4190 => x"80",
          4191 => x"82",
          4192 => x"91",
          4193 => x"90",
          4194 => x"82",
          4195 => x"85",
          4196 => x"9c",
          4197 => x"c2",
          4198 => x"0d",
          4199 => x"80",
          4200 => x"0b",
          4201 => x"84",
          4202 => x"b5",
          4203 => x"c0",
          4204 => x"04",
          4205 => x"76",
          4206 => x"98",
          4207 => x"2b",
          4208 => x"72",
          4209 => x"82",
          4210 => x"51",
          4211 => x"80",
          4212 => x"a8",
          4213 => x"53",
          4214 => x"9c",
          4215 => x"a4",
          4216 => x"02",
          4217 => x"05",
          4218 => x"52",
          4219 => x"72",
          4220 => x"06",
          4221 => x"53",
          4222 => x"98",
          4223 => x"0d",
          4224 => x"0d",
          4225 => x"05",
          4226 => x"71",
          4227 => x"54",
          4228 => x"b1",
          4229 => x"ec",
          4230 => x"51",
          4231 => x"3f",
          4232 => x"08",
          4233 => x"ff",
          4234 => x"82",
          4235 => x"52",
          4236 => x"ae",
          4237 => x"33",
          4238 => x"72",
          4239 => x"81",
          4240 => x"cc",
          4241 => x"ff",
          4242 => x"74",
          4243 => x"3d",
          4244 => x"3d",
          4245 => x"84",
          4246 => x"33",
          4247 => x"bb",
          4248 => x"b5",
          4249 => x"84",
          4250 => x"98",
          4251 => x"51",
          4252 => x"58",
          4253 => x"2e",
          4254 => x"51",
          4255 => x"82",
          4256 => x"70",
          4257 => x"b5",
          4258 => x"19",
          4259 => x"56",
          4260 => x"3f",
          4261 => x"08",
          4262 => x"b5",
          4263 => x"84",
          4264 => x"98",
          4265 => x"51",
          4266 => x"80",
          4267 => x"75",
          4268 => x"74",
          4269 => x"af",
          4270 => x"f0",
          4271 => x"55",
          4272 => x"f0",
          4273 => x"ff",
          4274 => x"75",
          4275 => x"80",
          4276 => x"f0",
          4277 => x"2e",
          4278 => x"b5",
          4279 => x"75",
          4280 => x"38",
          4281 => x"33",
          4282 => x"38",
          4283 => x"05",
          4284 => x"78",
          4285 => x"80",
          4286 => x"82",
          4287 => x"52",
          4288 => x"8f",
          4289 => x"b5",
          4290 => x"80",
          4291 => x"8c",
          4292 => x"fd",
          4293 => x"b5",
          4294 => x"54",
          4295 => x"71",
          4296 => x"38",
          4297 => x"d0",
          4298 => x"0c",
          4299 => x"14",
          4300 => x"80",
          4301 => x"80",
          4302 => x"f0",
          4303 => x"ec",
          4304 => x"80",
          4305 => x"71",
          4306 => x"c5",
          4307 => x"ec",
          4308 => x"a4",
          4309 => x"82",
          4310 => x"85",
          4311 => x"dc",
          4312 => x"57",
          4313 => x"b5",
          4314 => x"80",
          4315 => x"82",
          4316 => x"80",
          4317 => x"b5",
          4318 => x"80",
          4319 => x"3d",
          4320 => x"81",
          4321 => x"82",
          4322 => x"80",
          4323 => x"75",
          4324 => x"f3",
          4325 => x"98",
          4326 => x"0b",
          4327 => x"08",
          4328 => x"82",
          4329 => x"ff",
          4330 => x"55",
          4331 => x"34",
          4332 => x"52",
          4333 => x"ae",
          4334 => x"ff",
          4335 => x"74",
          4336 => x"81",
          4337 => x"38",
          4338 => x"04",
          4339 => x"aa",
          4340 => x"3d",
          4341 => x"81",
          4342 => x"80",
          4343 => x"ec",
          4344 => x"e2",
          4345 => x"b6",
          4346 => x"95",
          4347 => x"82",
          4348 => x"54",
          4349 => x"52",
          4350 => x"52",
          4351 => x"86",
          4352 => x"98",
          4353 => x"a5",
          4354 => x"ff",
          4355 => x"82",
          4356 => x"81",
          4357 => x"80",
          4358 => x"98",
          4359 => x"38",
          4360 => x"08",
          4361 => x"17",
          4362 => x"74",
          4363 => x"70",
          4364 => x"07",
          4365 => x"55",
          4366 => x"2e",
          4367 => x"ff",
          4368 => x"b5",
          4369 => x"11",
          4370 => x"80",
          4371 => x"82",
          4372 => x"80",
          4373 => x"82",
          4374 => x"ff",
          4375 => x"78",
          4376 => x"81",
          4377 => x"75",
          4378 => x"ff",
          4379 => x"79",
          4380 => x"93",
          4381 => x"08",
          4382 => x"98",
          4383 => x"80",
          4384 => x"b6",
          4385 => x"3d",
          4386 => x"3d",
          4387 => x"71",
          4388 => x"33",
          4389 => x"58",
          4390 => x"09",
          4391 => x"38",
          4392 => x"05",
          4393 => x"27",
          4394 => x"17",
          4395 => x"71",
          4396 => x"55",
          4397 => x"09",
          4398 => x"38",
          4399 => x"ea",
          4400 => x"73",
          4401 => x"b5",
          4402 => x"08",
          4403 => x"b2",
          4404 => x"b6",
          4405 => x"79",
          4406 => x"51",
          4407 => x"3f",
          4408 => x"08",
          4409 => x"84",
          4410 => x"74",
          4411 => x"38",
          4412 => x"88",
          4413 => x"fc",
          4414 => x"39",
          4415 => x"8c",
          4416 => x"53",
          4417 => x"c5",
          4418 => x"b6",
          4419 => x"2e",
          4420 => x"1b",
          4421 => x"77",
          4422 => x"3f",
          4423 => x"08",
          4424 => x"55",
          4425 => x"74",
          4426 => x"81",
          4427 => x"ff",
          4428 => x"82",
          4429 => x"8b",
          4430 => x"73",
          4431 => x"0c",
          4432 => x"04",
          4433 => x"b0",
          4434 => x"3d",
          4435 => x"08",
          4436 => x"80",
          4437 => x"34",
          4438 => x"33",
          4439 => x"08",
          4440 => x"81",
          4441 => x"82",
          4442 => x"55",
          4443 => x"38",
          4444 => x"80",
          4445 => x"38",
          4446 => x"06",
          4447 => x"80",
          4448 => x"38",
          4449 => x"86",
          4450 => x"98",
          4451 => x"ec",
          4452 => x"98",
          4453 => x"81",
          4454 => x"53",
          4455 => x"b6",
          4456 => x"80",
          4457 => x"82",
          4458 => x"80",
          4459 => x"82",
          4460 => x"ff",
          4461 => x"80",
          4462 => x"b6",
          4463 => x"82",
          4464 => x"53",
          4465 => x"90",
          4466 => x"54",
          4467 => x"3f",
          4468 => x"08",
          4469 => x"98",
          4470 => x"09",
          4471 => x"d0",
          4472 => x"98",
          4473 => x"b0",
          4474 => x"b6",
          4475 => x"80",
          4476 => x"98",
          4477 => x"38",
          4478 => x"08",
          4479 => x"17",
          4480 => x"74",
          4481 => x"74",
          4482 => x"52",
          4483 => x"c2",
          4484 => x"70",
          4485 => x"5c",
          4486 => x"27",
          4487 => x"5b",
          4488 => x"09",
          4489 => x"97",
          4490 => x"75",
          4491 => x"34",
          4492 => x"82",
          4493 => x"80",
          4494 => x"f9",
          4495 => x"3d",
          4496 => x"3f",
          4497 => x"08",
          4498 => x"98",
          4499 => x"78",
          4500 => x"38",
          4501 => x"06",
          4502 => x"33",
          4503 => x"70",
          4504 => x"cd",
          4505 => x"98",
          4506 => x"2c",
          4507 => x"05",
          4508 => x"82",
          4509 => x"70",
          4510 => x"33",
          4511 => x"51",
          4512 => x"59",
          4513 => x"56",
          4514 => x"80",
          4515 => x"74",
          4516 => x"74",
          4517 => x"29",
          4518 => x"05",
          4519 => x"51",
          4520 => x"24",
          4521 => x"76",
          4522 => x"77",
          4523 => x"3f",
          4524 => x"08",
          4525 => x"54",
          4526 => x"d7",
          4527 => x"cd",
          4528 => x"56",
          4529 => x"81",
          4530 => x"81",
          4531 => x"70",
          4532 => x"81",
          4533 => x"51",
          4534 => x"26",
          4535 => x"53",
          4536 => x"51",
          4537 => x"82",
          4538 => x"81",
          4539 => x"73",
          4540 => x"39",
          4541 => x"80",
          4542 => x"38",
          4543 => x"74",
          4544 => x"34",
          4545 => x"70",
          4546 => x"cd",
          4547 => x"98",
          4548 => x"2c",
          4549 => x"70",
          4550 => x"ab",
          4551 => x"5e",
          4552 => x"57",
          4553 => x"74",
          4554 => x"81",
          4555 => x"38",
          4556 => x"14",
          4557 => x"80",
          4558 => x"c4",
          4559 => x"82",
          4560 => x"92",
          4561 => x"cd",
          4562 => x"82",
          4563 => x"78",
          4564 => x"75",
          4565 => x"54",
          4566 => x"fd",
          4567 => x"84",
          4568 => x"b0",
          4569 => x"08",
          4570 => x"cc",
          4571 => x"7e",
          4572 => x"38",
          4573 => x"33",
          4574 => x"27",
          4575 => x"98",
          4576 => x"2c",
          4577 => x"75",
          4578 => x"74",
          4579 => x"33",
          4580 => x"74",
          4581 => x"29",
          4582 => x"05",
          4583 => x"82",
          4584 => x"56",
          4585 => x"39",
          4586 => x"33",
          4587 => x"54",
          4588 => x"cc",
          4589 => x"54",
          4590 => x"74",
          4591 => x"c8",
          4592 => x"7e",
          4593 => x"81",
          4594 => x"82",
          4595 => x"82",
          4596 => x"70",
          4597 => x"29",
          4598 => x"05",
          4599 => x"82",
          4600 => x"5a",
          4601 => x"74",
          4602 => x"38",
          4603 => x"08",
          4604 => x"70",
          4605 => x"ff",
          4606 => x"74",
          4607 => x"29",
          4608 => x"05",
          4609 => x"82",
          4610 => x"56",
          4611 => x"75",
          4612 => x"82",
          4613 => x"70",
          4614 => x"98",
          4615 => x"c8",
          4616 => x"56",
          4617 => x"25",
          4618 => x"82",
          4619 => x"52",
          4620 => x"a2",
          4621 => x"81",
          4622 => x"81",
          4623 => x"70",
          4624 => x"cd",
          4625 => x"51",
          4626 => x"24",
          4627 => x"ee",
          4628 => x"34",
          4629 => x"1b",
          4630 => x"cc",
          4631 => x"82",
          4632 => x"f3",
          4633 => x"fd",
          4634 => x"cc",
          4635 => x"ff",
          4636 => x"73",
          4637 => x"c6",
          4638 => x"c8",
          4639 => x"54",
          4640 => x"c8",
          4641 => x"54",
          4642 => x"cc",
          4643 => x"ec",
          4644 => x"51",
          4645 => x"3f",
          4646 => x"33",
          4647 => x"70",
          4648 => x"cd",
          4649 => x"51",
          4650 => x"74",
          4651 => x"74",
          4652 => x"14",
          4653 => x"82",
          4654 => x"52",
          4655 => x"ff",
          4656 => x"74",
          4657 => x"29",
          4658 => x"05",
          4659 => x"82",
          4660 => x"58",
          4661 => x"75",
          4662 => x"82",
          4663 => x"52",
          4664 => x"a1",
          4665 => x"cd",
          4666 => x"98",
          4667 => x"2c",
          4668 => x"33",
          4669 => x"57",
          4670 => x"fa",
          4671 => x"cd",
          4672 => x"88",
          4673 => x"ac",
          4674 => x"80",
          4675 => x"80",
          4676 => x"98",
          4677 => x"c8",
          4678 => x"55",
          4679 => x"de",
          4680 => x"39",
          4681 => x"33",
          4682 => x"80",
          4683 => x"cd",
          4684 => x"8a",
          4685 => x"fc",
          4686 => x"c8",
          4687 => x"f6",
          4688 => x"b6",
          4689 => x"ff",
          4690 => x"96",
          4691 => x"c8",
          4692 => x"80",
          4693 => x"81",
          4694 => x"79",
          4695 => x"3f",
          4696 => x"7a",
          4697 => x"82",
          4698 => x"80",
          4699 => x"c8",
          4700 => x"b6",
          4701 => x"3d",
          4702 => x"cd",
          4703 => x"73",
          4704 => x"ba",
          4705 => x"ec",
          4706 => x"51",
          4707 => x"3f",
          4708 => x"33",
          4709 => x"73",
          4710 => x"34",
          4711 => x"06",
          4712 => x"82",
          4713 => x"82",
          4714 => x"55",
          4715 => x"2e",
          4716 => x"ff",
          4717 => x"82",
          4718 => x"74",
          4719 => x"98",
          4720 => x"ff",
          4721 => x"55",
          4722 => x"ad",
          4723 => x"54",
          4724 => x"74",
          4725 => x"ec",
          4726 => x"33",
          4727 => x"d4",
          4728 => x"80",
          4729 => x"80",
          4730 => x"98",
          4731 => x"c8",
          4732 => x"55",
          4733 => x"d5",
          4734 => x"ec",
          4735 => x"51",
          4736 => x"3f",
          4737 => x"33",
          4738 => x"70",
          4739 => x"cd",
          4740 => x"51",
          4741 => x"74",
          4742 => x"38",
          4743 => x"08",
          4744 => x"ff",
          4745 => x"74",
          4746 => x"29",
          4747 => x"05",
          4748 => x"82",
          4749 => x"58",
          4750 => x"75",
          4751 => x"f7",
          4752 => x"cd",
          4753 => x"81",
          4754 => x"cd",
          4755 => x"56",
          4756 => x"27",
          4757 => x"82",
          4758 => x"52",
          4759 => x"73",
          4760 => x"34",
          4761 => x"33",
          4762 => x"9e",
          4763 => x"cd",
          4764 => x"81",
          4765 => x"cd",
          4766 => x"56",
          4767 => x"26",
          4768 => x"ba",
          4769 => x"cc",
          4770 => x"82",
          4771 => x"ee",
          4772 => x"0b",
          4773 => x"34",
          4774 => x"cd",
          4775 => x"9e",
          4776 => x"38",
          4777 => x"08",
          4778 => x"2e",
          4779 => x"51",
          4780 => x"3f",
          4781 => x"08",
          4782 => x"34",
          4783 => x"08",
          4784 => x"81",
          4785 => x"52",
          4786 => x"a8",
          4787 => x"5b",
          4788 => x"7a",
          4789 => x"b5",
          4790 => x"11",
          4791 => x"74",
          4792 => x"38",
          4793 => x"a6",
          4794 => x"b6",
          4795 => x"cd",
          4796 => x"b6",
          4797 => x"ff",
          4798 => x"53",
          4799 => x"51",
          4800 => x"3f",
          4801 => x"80",
          4802 => x"08",
          4803 => x"2e",
          4804 => x"74",
          4805 => x"ef",
          4806 => x"7a",
          4807 => x"81",
          4808 => x"82",
          4809 => x"55",
          4810 => x"a4",
          4811 => x"ff",
          4812 => x"82",
          4813 => x"82",
          4814 => x"82",
          4815 => x"81",
          4816 => x"05",
          4817 => x"79",
          4818 => x"9b",
          4819 => x"39",
          4820 => x"82",
          4821 => x"70",
          4822 => x"74",
          4823 => x"38",
          4824 => x"a5",
          4825 => x"b6",
          4826 => x"cd",
          4827 => x"b6",
          4828 => x"ff",
          4829 => x"53",
          4830 => x"51",
          4831 => x"3f",
          4832 => x"73",
          4833 => x"5b",
          4834 => x"82",
          4835 => x"74",
          4836 => x"cd",
          4837 => x"cd",
          4838 => x"79",
          4839 => x"3f",
          4840 => x"82",
          4841 => x"70",
          4842 => x"82",
          4843 => x"59",
          4844 => x"77",
          4845 => x"38",
          4846 => x"08",
          4847 => x"54",
          4848 => x"cc",
          4849 => x"70",
          4850 => x"ff",
          4851 => x"f4",
          4852 => x"cd",
          4853 => x"73",
          4854 => x"e2",
          4855 => x"ec",
          4856 => x"51",
          4857 => x"3f",
          4858 => x"33",
          4859 => x"73",
          4860 => x"34",
          4861 => x"f9",
          4862 => x"bf",
          4863 => x"b6",
          4864 => x"80",
          4865 => x"8c",
          4866 => x"53",
          4867 => x"bf",
          4868 => x"aa",
          4869 => x"b6",
          4870 => x"80",
          4871 => x"34",
          4872 => x"81",
          4873 => x"b6",
          4874 => x"77",
          4875 => x"76",
          4876 => x"82",
          4877 => x"54",
          4878 => x"34",
          4879 => x"34",
          4880 => x"08",
          4881 => x"22",
          4882 => x"80",
          4883 => x"83",
          4884 => x"70",
          4885 => x"51",
          4886 => x"88",
          4887 => x"89",
          4888 => x"b6",
          4889 => x"88",
          4890 => x"90",
          4891 => x"11",
          4892 => x"77",
          4893 => x"76",
          4894 => x"89",
          4895 => x"ff",
          4896 => x"52",
          4897 => x"72",
          4898 => x"fb",
          4899 => x"82",
          4900 => x"ff",
          4901 => x"51",
          4902 => x"b6",
          4903 => x"3d",
          4904 => x"3d",
          4905 => x"05",
          4906 => x"05",
          4907 => x"71",
          4908 => x"90",
          4909 => x"2b",
          4910 => x"83",
          4911 => x"70",
          4912 => x"33",
          4913 => x"07",
          4914 => x"ae",
          4915 => x"81",
          4916 => x"07",
          4917 => x"53",
          4918 => x"54",
          4919 => x"53",
          4920 => x"77",
          4921 => x"18",
          4922 => x"90",
          4923 => x"88",
          4924 => x"70",
          4925 => x"74",
          4926 => x"82",
          4927 => x"70",
          4928 => x"81",
          4929 => x"88",
          4930 => x"83",
          4931 => x"f8",
          4932 => x"56",
          4933 => x"73",
          4934 => x"06",
          4935 => x"54",
          4936 => x"82",
          4937 => x"81",
          4938 => x"72",
          4939 => x"82",
          4940 => x"16",
          4941 => x"34",
          4942 => x"34",
          4943 => x"04",
          4944 => x"82",
          4945 => x"02",
          4946 => x"05",
          4947 => x"2b",
          4948 => x"11",
          4949 => x"33",
          4950 => x"71",
          4951 => x"58",
          4952 => x"55",
          4953 => x"84",
          4954 => x"13",
          4955 => x"2b",
          4956 => x"2a",
          4957 => x"52",
          4958 => x"34",
          4959 => x"34",
          4960 => x"08",
          4961 => x"11",
          4962 => x"33",
          4963 => x"71",
          4964 => x"56",
          4965 => x"72",
          4966 => x"33",
          4967 => x"71",
          4968 => x"70",
          4969 => x"56",
          4970 => x"86",
          4971 => x"87",
          4972 => x"b6",
          4973 => x"70",
          4974 => x"33",
          4975 => x"07",
          4976 => x"ff",
          4977 => x"2a",
          4978 => x"53",
          4979 => x"34",
          4980 => x"34",
          4981 => x"04",
          4982 => x"02",
          4983 => x"82",
          4984 => x"71",
          4985 => x"11",
          4986 => x"12",
          4987 => x"2b",
          4988 => x"29",
          4989 => x"81",
          4990 => x"98",
          4991 => x"2b",
          4992 => x"53",
          4993 => x"56",
          4994 => x"71",
          4995 => x"f6",
          4996 => x"fe",
          4997 => x"b6",
          4998 => x"16",
          4999 => x"12",
          5000 => x"2b",
          5001 => x"07",
          5002 => x"33",
          5003 => x"71",
          5004 => x"70",
          5005 => x"ff",
          5006 => x"52",
          5007 => x"5a",
          5008 => x"05",
          5009 => x"54",
          5010 => x"13",
          5011 => x"13",
          5012 => x"90",
          5013 => x"70",
          5014 => x"33",
          5015 => x"71",
          5016 => x"56",
          5017 => x"72",
          5018 => x"81",
          5019 => x"88",
          5020 => x"81",
          5021 => x"70",
          5022 => x"51",
          5023 => x"72",
          5024 => x"81",
          5025 => x"3d",
          5026 => x"3d",
          5027 => x"90",
          5028 => x"05",
          5029 => x"70",
          5030 => x"11",
          5031 => x"83",
          5032 => x"8b",
          5033 => x"2b",
          5034 => x"59",
          5035 => x"73",
          5036 => x"81",
          5037 => x"88",
          5038 => x"8c",
          5039 => x"22",
          5040 => x"88",
          5041 => x"53",
          5042 => x"73",
          5043 => x"14",
          5044 => x"90",
          5045 => x"70",
          5046 => x"33",
          5047 => x"71",
          5048 => x"56",
          5049 => x"72",
          5050 => x"33",
          5051 => x"71",
          5052 => x"70",
          5053 => x"55",
          5054 => x"82",
          5055 => x"83",
          5056 => x"b6",
          5057 => x"82",
          5058 => x"12",
          5059 => x"2b",
          5060 => x"98",
          5061 => x"87",
          5062 => x"f7",
          5063 => x"82",
          5064 => x"31",
          5065 => x"83",
          5066 => x"70",
          5067 => x"fd",
          5068 => x"b6",
          5069 => x"83",
          5070 => x"82",
          5071 => x"12",
          5072 => x"2b",
          5073 => x"07",
          5074 => x"33",
          5075 => x"71",
          5076 => x"90",
          5077 => x"42",
          5078 => x"5b",
          5079 => x"54",
          5080 => x"8d",
          5081 => x"80",
          5082 => x"fe",
          5083 => x"84",
          5084 => x"33",
          5085 => x"71",
          5086 => x"83",
          5087 => x"11",
          5088 => x"53",
          5089 => x"55",
          5090 => x"34",
          5091 => x"06",
          5092 => x"14",
          5093 => x"90",
          5094 => x"84",
          5095 => x"13",
          5096 => x"2b",
          5097 => x"2a",
          5098 => x"56",
          5099 => x"16",
          5100 => x"16",
          5101 => x"90",
          5102 => x"80",
          5103 => x"34",
          5104 => x"14",
          5105 => x"90",
          5106 => x"84",
          5107 => x"85",
          5108 => x"b6",
          5109 => x"70",
          5110 => x"33",
          5111 => x"07",
          5112 => x"80",
          5113 => x"2a",
          5114 => x"56",
          5115 => x"34",
          5116 => x"34",
          5117 => x"04",
          5118 => x"73",
          5119 => x"90",
          5120 => x"f7",
          5121 => x"80",
          5122 => x"71",
          5123 => x"3f",
          5124 => x"04",
          5125 => x"80",
          5126 => x"f8",
          5127 => x"b6",
          5128 => x"ff",
          5129 => x"b6",
          5130 => x"11",
          5131 => x"33",
          5132 => x"07",
          5133 => x"56",
          5134 => x"ff",
          5135 => x"78",
          5136 => x"38",
          5137 => x"17",
          5138 => x"12",
          5139 => x"2b",
          5140 => x"ff",
          5141 => x"31",
          5142 => x"ff",
          5143 => x"27",
          5144 => x"56",
          5145 => x"79",
          5146 => x"73",
          5147 => x"38",
          5148 => x"5b",
          5149 => x"85",
          5150 => x"88",
          5151 => x"54",
          5152 => x"78",
          5153 => x"2e",
          5154 => x"79",
          5155 => x"76",
          5156 => x"b6",
          5157 => x"70",
          5158 => x"33",
          5159 => x"07",
          5160 => x"ff",
          5161 => x"5a",
          5162 => x"73",
          5163 => x"38",
          5164 => x"54",
          5165 => x"81",
          5166 => x"54",
          5167 => x"81",
          5168 => x"7a",
          5169 => x"06",
          5170 => x"51",
          5171 => x"81",
          5172 => x"80",
          5173 => x"52",
          5174 => x"c6",
          5175 => x"90",
          5176 => x"86",
          5177 => x"12",
          5178 => x"2b",
          5179 => x"07",
          5180 => x"55",
          5181 => x"17",
          5182 => x"ff",
          5183 => x"2a",
          5184 => x"54",
          5185 => x"34",
          5186 => x"06",
          5187 => x"15",
          5188 => x"90",
          5189 => x"2b",
          5190 => x"1e",
          5191 => x"87",
          5192 => x"88",
          5193 => x"88",
          5194 => x"5e",
          5195 => x"54",
          5196 => x"34",
          5197 => x"34",
          5198 => x"08",
          5199 => x"11",
          5200 => x"33",
          5201 => x"71",
          5202 => x"53",
          5203 => x"74",
          5204 => x"86",
          5205 => x"87",
          5206 => x"b6",
          5207 => x"16",
          5208 => x"11",
          5209 => x"33",
          5210 => x"07",
          5211 => x"53",
          5212 => x"56",
          5213 => x"16",
          5214 => x"16",
          5215 => x"90",
          5216 => x"05",
          5217 => x"b6",
          5218 => x"3d",
          5219 => x"3d",
          5220 => x"82",
          5221 => x"84",
          5222 => x"3f",
          5223 => x"80",
          5224 => x"71",
          5225 => x"3f",
          5226 => x"08",
          5227 => x"b6",
          5228 => x"3d",
          5229 => x"3d",
          5230 => x"40",
          5231 => x"42",
          5232 => x"90",
          5233 => x"09",
          5234 => x"38",
          5235 => x"7b",
          5236 => x"51",
          5237 => x"82",
          5238 => x"54",
          5239 => x"7e",
          5240 => x"51",
          5241 => x"7e",
          5242 => x"39",
          5243 => x"8f",
          5244 => x"98",
          5245 => x"ff",
          5246 => x"90",
          5247 => x"31",
          5248 => x"83",
          5249 => x"70",
          5250 => x"11",
          5251 => x"12",
          5252 => x"2b",
          5253 => x"31",
          5254 => x"ff",
          5255 => x"29",
          5256 => x"88",
          5257 => x"33",
          5258 => x"71",
          5259 => x"70",
          5260 => x"44",
          5261 => x"41",
          5262 => x"5b",
          5263 => x"5b",
          5264 => x"25",
          5265 => x"81",
          5266 => x"75",
          5267 => x"ff",
          5268 => x"54",
          5269 => x"83",
          5270 => x"88",
          5271 => x"88",
          5272 => x"33",
          5273 => x"71",
          5274 => x"90",
          5275 => x"47",
          5276 => x"54",
          5277 => x"8b",
          5278 => x"31",
          5279 => x"ff",
          5280 => x"77",
          5281 => x"fe",
          5282 => x"54",
          5283 => x"09",
          5284 => x"38",
          5285 => x"c0",
          5286 => x"ff",
          5287 => x"81",
          5288 => x"8e",
          5289 => x"24",
          5290 => x"51",
          5291 => x"81",
          5292 => x"18",
          5293 => x"24",
          5294 => x"79",
          5295 => x"33",
          5296 => x"71",
          5297 => x"53",
          5298 => x"f4",
          5299 => x"78",
          5300 => x"3f",
          5301 => x"08",
          5302 => x"06",
          5303 => x"53",
          5304 => x"82",
          5305 => x"11",
          5306 => x"55",
          5307 => x"ad",
          5308 => x"90",
          5309 => x"05",
          5310 => x"ff",
          5311 => x"81",
          5312 => x"15",
          5313 => x"24",
          5314 => x"78",
          5315 => x"3f",
          5316 => x"08",
          5317 => x"33",
          5318 => x"71",
          5319 => x"53",
          5320 => x"9c",
          5321 => x"78",
          5322 => x"3f",
          5323 => x"08",
          5324 => x"06",
          5325 => x"53",
          5326 => x"82",
          5327 => x"11",
          5328 => x"55",
          5329 => x"d5",
          5330 => x"90",
          5331 => x"05",
          5332 => x"19",
          5333 => x"83",
          5334 => x"58",
          5335 => x"7f",
          5336 => x"b0",
          5337 => x"98",
          5338 => x"b6",
          5339 => x"2e",
          5340 => x"53",
          5341 => x"b6",
          5342 => x"ff",
          5343 => x"73",
          5344 => x"3f",
          5345 => x"78",
          5346 => x"80",
          5347 => x"78",
          5348 => x"3f",
          5349 => x"2b",
          5350 => x"08",
          5351 => x"51",
          5352 => x"7b",
          5353 => x"b6",
          5354 => x"3d",
          5355 => x"3d",
          5356 => x"29",
          5357 => x"fb",
          5358 => x"b6",
          5359 => x"82",
          5360 => x"80",
          5361 => x"73",
          5362 => x"82",
          5363 => x"51",
          5364 => x"3f",
          5365 => x"98",
          5366 => x"0d",
          5367 => x"0d",
          5368 => x"33",
          5369 => x"70",
          5370 => x"38",
          5371 => x"11",
          5372 => x"82",
          5373 => x"83",
          5374 => x"fc",
          5375 => x"9b",
          5376 => x"84",
          5377 => x"33",
          5378 => x"51",
          5379 => x"80",
          5380 => x"84",
          5381 => x"92",
          5382 => x"51",
          5383 => x"80",
          5384 => x"81",
          5385 => x"72",
          5386 => x"92",
          5387 => x"81",
          5388 => x"0b",
          5389 => x"8c",
          5390 => x"71",
          5391 => x"06",
          5392 => x"80",
          5393 => x"87",
          5394 => x"08",
          5395 => x"38",
          5396 => x"80",
          5397 => x"71",
          5398 => x"c0",
          5399 => x"51",
          5400 => x"87",
          5401 => x"b6",
          5402 => x"82",
          5403 => x"33",
          5404 => x"b6",
          5405 => x"3d",
          5406 => x"3d",
          5407 => x"64",
          5408 => x"bf",
          5409 => x"40",
          5410 => x"74",
          5411 => x"cd",
          5412 => x"98",
          5413 => x"7a",
          5414 => x"81",
          5415 => x"72",
          5416 => x"87",
          5417 => x"11",
          5418 => x"8c",
          5419 => x"92",
          5420 => x"5a",
          5421 => x"58",
          5422 => x"c0",
          5423 => x"76",
          5424 => x"76",
          5425 => x"70",
          5426 => x"81",
          5427 => x"54",
          5428 => x"8e",
          5429 => x"52",
          5430 => x"81",
          5431 => x"81",
          5432 => x"74",
          5433 => x"53",
          5434 => x"83",
          5435 => x"78",
          5436 => x"8f",
          5437 => x"2e",
          5438 => x"c0",
          5439 => x"52",
          5440 => x"87",
          5441 => x"08",
          5442 => x"2e",
          5443 => x"84",
          5444 => x"38",
          5445 => x"87",
          5446 => x"15",
          5447 => x"70",
          5448 => x"52",
          5449 => x"ff",
          5450 => x"39",
          5451 => x"81",
          5452 => x"ff",
          5453 => x"57",
          5454 => x"90",
          5455 => x"80",
          5456 => x"71",
          5457 => x"78",
          5458 => x"38",
          5459 => x"80",
          5460 => x"80",
          5461 => x"81",
          5462 => x"72",
          5463 => x"0c",
          5464 => x"04",
          5465 => x"60",
          5466 => x"8c",
          5467 => x"33",
          5468 => x"5b",
          5469 => x"74",
          5470 => x"e1",
          5471 => x"98",
          5472 => x"79",
          5473 => x"78",
          5474 => x"06",
          5475 => x"77",
          5476 => x"87",
          5477 => x"11",
          5478 => x"8c",
          5479 => x"92",
          5480 => x"59",
          5481 => x"85",
          5482 => x"98",
          5483 => x"7d",
          5484 => x"0c",
          5485 => x"08",
          5486 => x"70",
          5487 => x"53",
          5488 => x"2e",
          5489 => x"70",
          5490 => x"33",
          5491 => x"18",
          5492 => x"2a",
          5493 => x"51",
          5494 => x"2e",
          5495 => x"c0",
          5496 => x"52",
          5497 => x"87",
          5498 => x"08",
          5499 => x"2e",
          5500 => x"84",
          5501 => x"38",
          5502 => x"87",
          5503 => x"15",
          5504 => x"70",
          5505 => x"52",
          5506 => x"ff",
          5507 => x"39",
          5508 => x"81",
          5509 => x"80",
          5510 => x"52",
          5511 => x"90",
          5512 => x"80",
          5513 => x"71",
          5514 => x"7a",
          5515 => x"38",
          5516 => x"80",
          5517 => x"80",
          5518 => x"81",
          5519 => x"72",
          5520 => x"0c",
          5521 => x"04",
          5522 => x"7a",
          5523 => x"a3",
          5524 => x"88",
          5525 => x"33",
          5526 => x"56",
          5527 => x"3f",
          5528 => x"08",
          5529 => x"83",
          5530 => x"fe",
          5531 => x"87",
          5532 => x"0c",
          5533 => x"76",
          5534 => x"38",
          5535 => x"93",
          5536 => x"2b",
          5537 => x"8c",
          5538 => x"71",
          5539 => x"38",
          5540 => x"71",
          5541 => x"c6",
          5542 => x"39",
          5543 => x"81",
          5544 => x"06",
          5545 => x"71",
          5546 => x"38",
          5547 => x"8c",
          5548 => x"e8",
          5549 => x"98",
          5550 => x"71",
          5551 => x"73",
          5552 => x"92",
          5553 => x"72",
          5554 => x"06",
          5555 => x"f7",
          5556 => x"80",
          5557 => x"88",
          5558 => x"0c",
          5559 => x"80",
          5560 => x"56",
          5561 => x"56",
          5562 => x"82",
          5563 => x"88",
          5564 => x"fe",
          5565 => x"81",
          5566 => x"33",
          5567 => x"07",
          5568 => x"0c",
          5569 => x"3d",
          5570 => x"3d",
          5571 => x"11",
          5572 => x"33",
          5573 => x"71",
          5574 => x"81",
          5575 => x"72",
          5576 => x"75",
          5577 => x"82",
          5578 => x"52",
          5579 => x"54",
          5580 => x"0d",
          5581 => x"0d",
          5582 => x"05",
          5583 => x"52",
          5584 => x"70",
          5585 => x"34",
          5586 => x"51",
          5587 => x"83",
          5588 => x"ff",
          5589 => x"75",
          5590 => x"72",
          5591 => x"54",
          5592 => x"2a",
          5593 => x"70",
          5594 => x"34",
          5595 => x"51",
          5596 => x"81",
          5597 => x"70",
          5598 => x"70",
          5599 => x"3d",
          5600 => x"3d",
          5601 => x"77",
          5602 => x"70",
          5603 => x"38",
          5604 => x"05",
          5605 => x"70",
          5606 => x"34",
          5607 => x"eb",
          5608 => x"0d",
          5609 => x"0d",
          5610 => x"54",
          5611 => x"72",
          5612 => x"54",
          5613 => x"51",
          5614 => x"84",
          5615 => x"fc",
          5616 => x"77",
          5617 => x"53",
          5618 => x"05",
          5619 => x"70",
          5620 => x"33",
          5621 => x"ff",
          5622 => x"52",
          5623 => x"2e",
          5624 => x"80",
          5625 => x"71",
          5626 => x"0c",
          5627 => x"04",
          5628 => x"74",
          5629 => x"89",
          5630 => x"2e",
          5631 => x"11",
          5632 => x"52",
          5633 => x"70",
          5634 => x"98",
          5635 => x"0d",
          5636 => x"82",
          5637 => x"04",
          5638 => x"b6",
          5639 => x"f7",
          5640 => x"56",
          5641 => x"17",
          5642 => x"74",
          5643 => x"d6",
          5644 => x"b0",
          5645 => x"b4",
          5646 => x"81",
          5647 => x"59",
          5648 => x"82",
          5649 => x"7a",
          5650 => x"06",
          5651 => x"b6",
          5652 => x"17",
          5653 => x"08",
          5654 => x"08",
          5655 => x"08",
          5656 => x"74",
          5657 => x"38",
          5658 => x"55",
          5659 => x"09",
          5660 => x"38",
          5661 => x"18",
          5662 => x"81",
          5663 => x"f9",
          5664 => x"39",
          5665 => x"82",
          5666 => x"8b",
          5667 => x"fa",
          5668 => x"7a",
          5669 => x"57",
          5670 => x"08",
          5671 => x"75",
          5672 => x"3f",
          5673 => x"08",
          5674 => x"98",
          5675 => x"81",
          5676 => x"b4",
          5677 => x"16",
          5678 => x"be",
          5679 => x"98",
          5680 => x"85",
          5681 => x"81",
          5682 => x"17",
          5683 => x"b6",
          5684 => x"3d",
          5685 => x"3d",
          5686 => x"52",
          5687 => x"3f",
          5688 => x"08",
          5689 => x"98",
          5690 => x"38",
          5691 => x"74",
          5692 => x"81",
          5693 => x"38",
          5694 => x"59",
          5695 => x"09",
          5696 => x"e3",
          5697 => x"53",
          5698 => x"08",
          5699 => x"70",
          5700 => x"91",
          5701 => x"d5",
          5702 => x"17",
          5703 => x"3f",
          5704 => x"a4",
          5705 => x"51",
          5706 => x"86",
          5707 => x"f2",
          5708 => x"17",
          5709 => x"3f",
          5710 => x"52",
          5711 => x"51",
          5712 => x"8c",
          5713 => x"84",
          5714 => x"fc",
          5715 => x"17",
          5716 => x"70",
          5717 => x"79",
          5718 => x"52",
          5719 => x"51",
          5720 => x"77",
          5721 => x"80",
          5722 => x"81",
          5723 => x"f9",
          5724 => x"b6",
          5725 => x"2e",
          5726 => x"58",
          5727 => x"98",
          5728 => x"0d",
          5729 => x"0d",
          5730 => x"98",
          5731 => x"05",
          5732 => x"80",
          5733 => x"27",
          5734 => x"14",
          5735 => x"29",
          5736 => x"05",
          5737 => x"82",
          5738 => x"87",
          5739 => x"f9",
          5740 => x"7a",
          5741 => x"54",
          5742 => x"27",
          5743 => x"76",
          5744 => x"27",
          5745 => x"ff",
          5746 => x"58",
          5747 => x"80",
          5748 => x"82",
          5749 => x"72",
          5750 => x"38",
          5751 => x"72",
          5752 => x"8e",
          5753 => x"39",
          5754 => x"17",
          5755 => x"a4",
          5756 => x"53",
          5757 => x"fd",
          5758 => x"b6",
          5759 => x"9f",
          5760 => x"ff",
          5761 => x"11",
          5762 => x"70",
          5763 => x"18",
          5764 => x"76",
          5765 => x"53",
          5766 => x"82",
          5767 => x"80",
          5768 => x"83",
          5769 => x"b4",
          5770 => x"88",
          5771 => x"79",
          5772 => x"84",
          5773 => x"58",
          5774 => x"80",
          5775 => x"9f",
          5776 => x"80",
          5777 => x"88",
          5778 => x"08",
          5779 => x"51",
          5780 => x"82",
          5781 => x"80",
          5782 => x"10",
          5783 => x"74",
          5784 => x"51",
          5785 => x"82",
          5786 => x"83",
          5787 => x"58",
          5788 => x"87",
          5789 => x"08",
          5790 => x"51",
          5791 => x"82",
          5792 => x"9b",
          5793 => x"2b",
          5794 => x"74",
          5795 => x"51",
          5796 => x"82",
          5797 => x"f0",
          5798 => x"83",
          5799 => x"77",
          5800 => x"0c",
          5801 => x"04",
          5802 => x"7a",
          5803 => x"58",
          5804 => x"81",
          5805 => x"9e",
          5806 => x"17",
          5807 => x"96",
          5808 => x"53",
          5809 => x"81",
          5810 => x"79",
          5811 => x"72",
          5812 => x"38",
          5813 => x"72",
          5814 => x"b8",
          5815 => x"39",
          5816 => x"17",
          5817 => x"a4",
          5818 => x"53",
          5819 => x"fb",
          5820 => x"b6",
          5821 => x"82",
          5822 => x"81",
          5823 => x"83",
          5824 => x"b4",
          5825 => x"78",
          5826 => x"56",
          5827 => x"76",
          5828 => x"38",
          5829 => x"9f",
          5830 => x"33",
          5831 => x"07",
          5832 => x"74",
          5833 => x"83",
          5834 => x"89",
          5835 => x"08",
          5836 => x"51",
          5837 => x"82",
          5838 => x"59",
          5839 => x"08",
          5840 => x"74",
          5841 => x"16",
          5842 => x"84",
          5843 => x"76",
          5844 => x"88",
          5845 => x"81",
          5846 => x"8f",
          5847 => x"53",
          5848 => x"80",
          5849 => x"88",
          5850 => x"08",
          5851 => x"51",
          5852 => x"82",
          5853 => x"59",
          5854 => x"08",
          5855 => x"77",
          5856 => x"06",
          5857 => x"83",
          5858 => x"05",
          5859 => x"f7",
          5860 => x"39",
          5861 => x"a4",
          5862 => x"52",
          5863 => x"ef",
          5864 => x"98",
          5865 => x"b6",
          5866 => x"38",
          5867 => x"06",
          5868 => x"83",
          5869 => x"18",
          5870 => x"54",
          5871 => x"f6",
          5872 => x"b6",
          5873 => x"0a",
          5874 => x"52",
          5875 => x"83",
          5876 => x"83",
          5877 => x"82",
          5878 => x"8a",
          5879 => x"f8",
          5880 => x"7c",
          5881 => x"59",
          5882 => x"81",
          5883 => x"38",
          5884 => x"08",
          5885 => x"73",
          5886 => x"38",
          5887 => x"52",
          5888 => x"a4",
          5889 => x"98",
          5890 => x"b6",
          5891 => x"f2",
          5892 => x"82",
          5893 => x"39",
          5894 => x"e6",
          5895 => x"98",
          5896 => x"de",
          5897 => x"78",
          5898 => x"3f",
          5899 => x"08",
          5900 => x"98",
          5901 => x"80",
          5902 => x"b6",
          5903 => x"2e",
          5904 => x"b6",
          5905 => x"2e",
          5906 => x"53",
          5907 => x"51",
          5908 => x"82",
          5909 => x"c5",
          5910 => x"08",
          5911 => x"18",
          5912 => x"57",
          5913 => x"90",
          5914 => x"90",
          5915 => x"16",
          5916 => x"54",
          5917 => x"34",
          5918 => x"78",
          5919 => x"38",
          5920 => x"82",
          5921 => x"8a",
          5922 => x"f6",
          5923 => x"7e",
          5924 => x"5b",
          5925 => x"38",
          5926 => x"58",
          5927 => x"88",
          5928 => x"08",
          5929 => x"38",
          5930 => x"39",
          5931 => x"51",
          5932 => x"81",
          5933 => x"b6",
          5934 => x"82",
          5935 => x"b6",
          5936 => x"82",
          5937 => x"ff",
          5938 => x"38",
          5939 => x"82",
          5940 => x"26",
          5941 => x"79",
          5942 => x"08",
          5943 => x"73",
          5944 => x"b9",
          5945 => x"2e",
          5946 => x"80",
          5947 => x"1a",
          5948 => x"08",
          5949 => x"38",
          5950 => x"52",
          5951 => x"af",
          5952 => x"82",
          5953 => x"81",
          5954 => x"06",
          5955 => x"b6",
          5956 => x"82",
          5957 => x"09",
          5958 => x"72",
          5959 => x"70",
          5960 => x"b6",
          5961 => x"51",
          5962 => x"73",
          5963 => x"82",
          5964 => x"80",
          5965 => x"8c",
          5966 => x"81",
          5967 => x"38",
          5968 => x"08",
          5969 => x"73",
          5970 => x"75",
          5971 => x"77",
          5972 => x"56",
          5973 => x"76",
          5974 => x"82",
          5975 => x"26",
          5976 => x"75",
          5977 => x"f8",
          5978 => x"b6",
          5979 => x"2e",
          5980 => x"59",
          5981 => x"08",
          5982 => x"81",
          5983 => x"82",
          5984 => x"59",
          5985 => x"08",
          5986 => x"70",
          5987 => x"25",
          5988 => x"51",
          5989 => x"73",
          5990 => x"75",
          5991 => x"81",
          5992 => x"38",
          5993 => x"f5",
          5994 => x"75",
          5995 => x"f9",
          5996 => x"b6",
          5997 => x"b6",
          5998 => x"70",
          5999 => x"08",
          6000 => x"51",
          6001 => x"80",
          6002 => x"73",
          6003 => x"38",
          6004 => x"52",
          6005 => x"d0",
          6006 => x"98",
          6007 => x"a5",
          6008 => x"18",
          6009 => x"08",
          6010 => x"18",
          6011 => x"74",
          6012 => x"38",
          6013 => x"18",
          6014 => x"33",
          6015 => x"73",
          6016 => x"97",
          6017 => x"74",
          6018 => x"38",
          6019 => x"55",
          6020 => x"b6",
          6021 => x"85",
          6022 => x"75",
          6023 => x"b6",
          6024 => x"3d",
          6025 => x"3d",
          6026 => x"52",
          6027 => x"3f",
          6028 => x"08",
          6029 => x"82",
          6030 => x"80",
          6031 => x"52",
          6032 => x"c1",
          6033 => x"98",
          6034 => x"98",
          6035 => x"0c",
          6036 => x"53",
          6037 => x"15",
          6038 => x"f2",
          6039 => x"56",
          6040 => x"16",
          6041 => x"22",
          6042 => x"27",
          6043 => x"54",
          6044 => x"76",
          6045 => x"33",
          6046 => x"3f",
          6047 => x"08",
          6048 => x"38",
          6049 => x"76",
          6050 => x"70",
          6051 => x"9f",
          6052 => x"56",
          6053 => x"b6",
          6054 => x"3d",
          6055 => x"3d",
          6056 => x"71",
          6057 => x"57",
          6058 => x"0a",
          6059 => x"38",
          6060 => x"53",
          6061 => x"38",
          6062 => x"0c",
          6063 => x"54",
          6064 => x"75",
          6065 => x"73",
          6066 => x"a8",
          6067 => x"73",
          6068 => x"85",
          6069 => x"0b",
          6070 => x"5a",
          6071 => x"27",
          6072 => x"a8",
          6073 => x"18",
          6074 => x"39",
          6075 => x"70",
          6076 => x"58",
          6077 => x"b2",
          6078 => x"76",
          6079 => x"3f",
          6080 => x"08",
          6081 => x"98",
          6082 => x"bd",
          6083 => x"82",
          6084 => x"27",
          6085 => x"16",
          6086 => x"98",
          6087 => x"38",
          6088 => x"39",
          6089 => x"55",
          6090 => x"52",
          6091 => x"d5",
          6092 => x"98",
          6093 => x"0c",
          6094 => x"0c",
          6095 => x"53",
          6096 => x"80",
          6097 => x"85",
          6098 => x"94",
          6099 => x"2a",
          6100 => x"0c",
          6101 => x"06",
          6102 => x"9c",
          6103 => x"58",
          6104 => x"98",
          6105 => x"0d",
          6106 => x"0d",
          6107 => x"90",
          6108 => x"05",
          6109 => x"f0",
          6110 => x"27",
          6111 => x"0b",
          6112 => x"98",
          6113 => x"84",
          6114 => x"2e",
          6115 => x"76",
          6116 => x"58",
          6117 => x"38",
          6118 => x"15",
          6119 => x"08",
          6120 => x"38",
          6121 => x"88",
          6122 => x"53",
          6123 => x"81",
          6124 => x"c0",
          6125 => x"22",
          6126 => x"89",
          6127 => x"72",
          6128 => x"74",
          6129 => x"f3",
          6130 => x"b6",
          6131 => x"82",
          6132 => x"82",
          6133 => x"27",
          6134 => x"81",
          6135 => x"98",
          6136 => x"80",
          6137 => x"16",
          6138 => x"98",
          6139 => x"ca",
          6140 => x"38",
          6141 => x"0c",
          6142 => x"dd",
          6143 => x"08",
          6144 => x"f9",
          6145 => x"b6",
          6146 => x"87",
          6147 => x"98",
          6148 => x"80",
          6149 => x"55",
          6150 => x"08",
          6151 => x"38",
          6152 => x"b6",
          6153 => x"2e",
          6154 => x"b6",
          6155 => x"75",
          6156 => x"3f",
          6157 => x"08",
          6158 => x"94",
          6159 => x"52",
          6160 => x"c1",
          6161 => x"98",
          6162 => x"0c",
          6163 => x"0c",
          6164 => x"05",
          6165 => x"80",
          6166 => x"b6",
          6167 => x"3d",
          6168 => x"3d",
          6169 => x"71",
          6170 => x"57",
          6171 => x"51",
          6172 => x"82",
          6173 => x"54",
          6174 => x"08",
          6175 => x"82",
          6176 => x"56",
          6177 => x"52",
          6178 => x"83",
          6179 => x"98",
          6180 => x"b6",
          6181 => x"d2",
          6182 => x"98",
          6183 => x"08",
          6184 => x"54",
          6185 => x"e5",
          6186 => x"06",
          6187 => x"58",
          6188 => x"08",
          6189 => x"38",
          6190 => x"75",
          6191 => x"80",
          6192 => x"81",
          6193 => x"7a",
          6194 => x"06",
          6195 => x"39",
          6196 => x"08",
          6197 => x"76",
          6198 => x"3f",
          6199 => x"08",
          6200 => x"98",
          6201 => x"ff",
          6202 => x"84",
          6203 => x"06",
          6204 => x"54",
          6205 => x"98",
          6206 => x"0d",
          6207 => x"0d",
          6208 => x"52",
          6209 => x"3f",
          6210 => x"08",
          6211 => x"06",
          6212 => x"51",
          6213 => x"83",
          6214 => x"06",
          6215 => x"14",
          6216 => x"3f",
          6217 => x"08",
          6218 => x"07",
          6219 => x"b6",
          6220 => x"3d",
          6221 => x"3d",
          6222 => x"70",
          6223 => x"06",
          6224 => x"53",
          6225 => x"ed",
          6226 => x"33",
          6227 => x"83",
          6228 => x"06",
          6229 => x"90",
          6230 => x"15",
          6231 => x"3f",
          6232 => x"04",
          6233 => x"7b",
          6234 => x"84",
          6235 => x"58",
          6236 => x"80",
          6237 => x"38",
          6238 => x"52",
          6239 => x"8f",
          6240 => x"98",
          6241 => x"b6",
          6242 => x"f5",
          6243 => x"08",
          6244 => x"53",
          6245 => x"84",
          6246 => x"39",
          6247 => x"70",
          6248 => x"81",
          6249 => x"51",
          6250 => x"16",
          6251 => x"98",
          6252 => x"81",
          6253 => x"38",
          6254 => x"ae",
          6255 => x"81",
          6256 => x"54",
          6257 => x"2e",
          6258 => x"8f",
          6259 => x"82",
          6260 => x"76",
          6261 => x"54",
          6262 => x"09",
          6263 => x"38",
          6264 => x"7a",
          6265 => x"80",
          6266 => x"fa",
          6267 => x"b6",
          6268 => x"82",
          6269 => x"89",
          6270 => x"08",
          6271 => x"86",
          6272 => x"98",
          6273 => x"82",
          6274 => x"8b",
          6275 => x"fb",
          6276 => x"70",
          6277 => x"81",
          6278 => x"fc",
          6279 => x"b6",
          6280 => x"82",
          6281 => x"b4",
          6282 => x"08",
          6283 => x"ec",
          6284 => x"b6",
          6285 => x"82",
          6286 => x"a0",
          6287 => x"82",
          6288 => x"52",
          6289 => x"51",
          6290 => x"8b",
          6291 => x"52",
          6292 => x"51",
          6293 => x"81",
          6294 => x"34",
          6295 => x"98",
          6296 => x"0d",
          6297 => x"0d",
          6298 => x"98",
          6299 => x"70",
          6300 => x"ec",
          6301 => x"b6",
          6302 => x"38",
          6303 => x"53",
          6304 => x"81",
          6305 => x"34",
          6306 => x"04",
          6307 => x"78",
          6308 => x"80",
          6309 => x"34",
          6310 => x"80",
          6311 => x"38",
          6312 => x"18",
          6313 => x"9c",
          6314 => x"70",
          6315 => x"56",
          6316 => x"a0",
          6317 => x"71",
          6318 => x"81",
          6319 => x"81",
          6320 => x"89",
          6321 => x"06",
          6322 => x"73",
          6323 => x"55",
          6324 => x"55",
          6325 => x"81",
          6326 => x"81",
          6327 => x"74",
          6328 => x"75",
          6329 => x"52",
          6330 => x"13",
          6331 => x"08",
          6332 => x"33",
          6333 => x"9c",
          6334 => x"11",
          6335 => x"8a",
          6336 => x"98",
          6337 => x"96",
          6338 => x"e7",
          6339 => x"98",
          6340 => x"23",
          6341 => x"e7",
          6342 => x"b6",
          6343 => x"17",
          6344 => x"0d",
          6345 => x"0d",
          6346 => x"5e",
          6347 => x"70",
          6348 => x"55",
          6349 => x"83",
          6350 => x"73",
          6351 => x"91",
          6352 => x"2e",
          6353 => x"1d",
          6354 => x"0c",
          6355 => x"15",
          6356 => x"70",
          6357 => x"56",
          6358 => x"09",
          6359 => x"38",
          6360 => x"80",
          6361 => x"30",
          6362 => x"78",
          6363 => x"54",
          6364 => x"73",
          6365 => x"60",
          6366 => x"54",
          6367 => x"96",
          6368 => x"0b",
          6369 => x"80",
          6370 => x"f6",
          6371 => x"b6",
          6372 => x"85",
          6373 => x"3d",
          6374 => x"5c",
          6375 => x"53",
          6376 => x"51",
          6377 => x"80",
          6378 => x"88",
          6379 => x"5c",
          6380 => x"09",
          6381 => x"d4",
          6382 => x"70",
          6383 => x"71",
          6384 => x"30",
          6385 => x"73",
          6386 => x"51",
          6387 => x"57",
          6388 => x"38",
          6389 => x"75",
          6390 => x"17",
          6391 => x"75",
          6392 => x"30",
          6393 => x"51",
          6394 => x"80",
          6395 => x"38",
          6396 => x"87",
          6397 => x"26",
          6398 => x"77",
          6399 => x"a4",
          6400 => x"27",
          6401 => x"a0",
          6402 => x"39",
          6403 => x"33",
          6404 => x"57",
          6405 => x"27",
          6406 => x"75",
          6407 => x"30",
          6408 => x"32",
          6409 => x"80",
          6410 => x"25",
          6411 => x"56",
          6412 => x"80",
          6413 => x"84",
          6414 => x"58",
          6415 => x"70",
          6416 => x"55",
          6417 => x"09",
          6418 => x"38",
          6419 => x"80",
          6420 => x"30",
          6421 => x"77",
          6422 => x"54",
          6423 => x"81",
          6424 => x"ae",
          6425 => x"06",
          6426 => x"54",
          6427 => x"74",
          6428 => x"80",
          6429 => x"7b",
          6430 => x"30",
          6431 => x"70",
          6432 => x"25",
          6433 => x"07",
          6434 => x"51",
          6435 => x"a7",
          6436 => x"8b",
          6437 => x"39",
          6438 => x"54",
          6439 => x"8c",
          6440 => x"ff",
          6441 => x"e0",
          6442 => x"54",
          6443 => x"e1",
          6444 => x"98",
          6445 => x"b2",
          6446 => x"70",
          6447 => x"71",
          6448 => x"54",
          6449 => x"82",
          6450 => x"80",
          6451 => x"38",
          6452 => x"76",
          6453 => x"df",
          6454 => x"54",
          6455 => x"81",
          6456 => x"55",
          6457 => x"34",
          6458 => x"52",
          6459 => x"51",
          6460 => x"82",
          6461 => x"bf",
          6462 => x"16",
          6463 => x"26",
          6464 => x"16",
          6465 => x"06",
          6466 => x"17",
          6467 => x"34",
          6468 => x"fd",
          6469 => x"19",
          6470 => x"80",
          6471 => x"79",
          6472 => x"81",
          6473 => x"81",
          6474 => x"85",
          6475 => x"54",
          6476 => x"8f",
          6477 => x"86",
          6478 => x"39",
          6479 => x"f3",
          6480 => x"73",
          6481 => x"80",
          6482 => x"52",
          6483 => x"ce",
          6484 => x"98",
          6485 => x"b6",
          6486 => x"d7",
          6487 => x"08",
          6488 => x"e6",
          6489 => x"b6",
          6490 => x"82",
          6491 => x"80",
          6492 => x"1b",
          6493 => x"55",
          6494 => x"2e",
          6495 => x"8b",
          6496 => x"06",
          6497 => x"1c",
          6498 => x"33",
          6499 => x"70",
          6500 => x"55",
          6501 => x"38",
          6502 => x"52",
          6503 => x"9f",
          6504 => x"98",
          6505 => x"8b",
          6506 => x"7a",
          6507 => x"3f",
          6508 => x"75",
          6509 => x"57",
          6510 => x"2e",
          6511 => x"84",
          6512 => x"06",
          6513 => x"75",
          6514 => x"81",
          6515 => x"2a",
          6516 => x"73",
          6517 => x"38",
          6518 => x"54",
          6519 => x"fb",
          6520 => x"80",
          6521 => x"34",
          6522 => x"c1",
          6523 => x"06",
          6524 => x"38",
          6525 => x"39",
          6526 => x"70",
          6527 => x"54",
          6528 => x"86",
          6529 => x"84",
          6530 => x"06",
          6531 => x"73",
          6532 => x"38",
          6533 => x"83",
          6534 => x"b4",
          6535 => x"51",
          6536 => x"82",
          6537 => x"88",
          6538 => x"ea",
          6539 => x"b6",
          6540 => x"3d",
          6541 => x"3d",
          6542 => x"ff",
          6543 => x"71",
          6544 => x"5c",
          6545 => x"80",
          6546 => x"38",
          6547 => x"05",
          6548 => x"a0",
          6549 => x"71",
          6550 => x"38",
          6551 => x"71",
          6552 => x"81",
          6553 => x"38",
          6554 => x"11",
          6555 => x"06",
          6556 => x"70",
          6557 => x"38",
          6558 => x"81",
          6559 => x"05",
          6560 => x"76",
          6561 => x"38",
          6562 => x"af",
          6563 => x"77",
          6564 => x"57",
          6565 => x"05",
          6566 => x"70",
          6567 => x"33",
          6568 => x"53",
          6569 => x"99",
          6570 => x"e0",
          6571 => x"ff",
          6572 => x"ff",
          6573 => x"70",
          6574 => x"38",
          6575 => x"81",
          6576 => x"51",
          6577 => x"9f",
          6578 => x"72",
          6579 => x"81",
          6580 => x"70",
          6581 => x"72",
          6582 => x"32",
          6583 => x"72",
          6584 => x"73",
          6585 => x"53",
          6586 => x"70",
          6587 => x"38",
          6588 => x"19",
          6589 => x"75",
          6590 => x"38",
          6591 => x"83",
          6592 => x"74",
          6593 => x"59",
          6594 => x"39",
          6595 => x"33",
          6596 => x"b6",
          6597 => x"3d",
          6598 => x"3d",
          6599 => x"80",
          6600 => x"34",
          6601 => x"17",
          6602 => x"75",
          6603 => x"3f",
          6604 => x"b6",
          6605 => x"80",
          6606 => x"16",
          6607 => x"3f",
          6608 => x"08",
          6609 => x"06",
          6610 => x"73",
          6611 => x"2e",
          6612 => x"80",
          6613 => x"0b",
          6614 => x"56",
          6615 => x"e9",
          6616 => x"06",
          6617 => x"57",
          6618 => x"32",
          6619 => x"80",
          6620 => x"51",
          6621 => x"8a",
          6622 => x"e8",
          6623 => x"06",
          6624 => x"53",
          6625 => x"52",
          6626 => x"51",
          6627 => x"82",
          6628 => x"55",
          6629 => x"08",
          6630 => x"38",
          6631 => x"af",
          6632 => x"86",
          6633 => x"97",
          6634 => x"98",
          6635 => x"b6",
          6636 => x"2e",
          6637 => x"55",
          6638 => x"98",
          6639 => x"0d",
          6640 => x"0d",
          6641 => x"05",
          6642 => x"33",
          6643 => x"75",
          6644 => x"fc",
          6645 => x"b6",
          6646 => x"8b",
          6647 => x"82",
          6648 => x"24",
          6649 => x"82",
          6650 => x"84",
          6651 => x"d0",
          6652 => x"55",
          6653 => x"73",
          6654 => x"e6",
          6655 => x"0c",
          6656 => x"06",
          6657 => x"57",
          6658 => x"ae",
          6659 => x"33",
          6660 => x"3f",
          6661 => x"08",
          6662 => x"70",
          6663 => x"55",
          6664 => x"76",
          6665 => x"b8",
          6666 => x"2a",
          6667 => x"51",
          6668 => x"72",
          6669 => x"86",
          6670 => x"74",
          6671 => x"15",
          6672 => x"81",
          6673 => x"d7",
          6674 => x"b6",
          6675 => x"ff",
          6676 => x"06",
          6677 => x"56",
          6678 => x"38",
          6679 => x"8f",
          6680 => x"2a",
          6681 => x"51",
          6682 => x"72",
          6683 => x"80",
          6684 => x"52",
          6685 => x"3f",
          6686 => x"08",
          6687 => x"57",
          6688 => x"09",
          6689 => x"e2",
          6690 => x"74",
          6691 => x"56",
          6692 => x"33",
          6693 => x"72",
          6694 => x"38",
          6695 => x"51",
          6696 => x"82",
          6697 => x"57",
          6698 => x"84",
          6699 => x"ff",
          6700 => x"56",
          6701 => x"25",
          6702 => x"0b",
          6703 => x"56",
          6704 => x"05",
          6705 => x"83",
          6706 => x"2e",
          6707 => x"52",
          6708 => x"c6",
          6709 => x"98",
          6710 => x"06",
          6711 => x"27",
          6712 => x"16",
          6713 => x"27",
          6714 => x"56",
          6715 => x"84",
          6716 => x"56",
          6717 => x"84",
          6718 => x"14",
          6719 => x"3f",
          6720 => x"08",
          6721 => x"06",
          6722 => x"80",
          6723 => x"06",
          6724 => x"80",
          6725 => x"db",
          6726 => x"b6",
          6727 => x"ff",
          6728 => x"77",
          6729 => x"d8",
          6730 => x"de",
          6731 => x"98",
          6732 => x"9c",
          6733 => x"c4",
          6734 => x"15",
          6735 => x"14",
          6736 => x"70",
          6737 => x"51",
          6738 => x"56",
          6739 => x"84",
          6740 => x"81",
          6741 => x"71",
          6742 => x"16",
          6743 => x"53",
          6744 => x"23",
          6745 => x"8b",
          6746 => x"73",
          6747 => x"80",
          6748 => x"8d",
          6749 => x"39",
          6750 => x"51",
          6751 => x"82",
          6752 => x"53",
          6753 => x"08",
          6754 => x"72",
          6755 => x"8d",
          6756 => x"ce",
          6757 => x"14",
          6758 => x"3f",
          6759 => x"08",
          6760 => x"06",
          6761 => x"38",
          6762 => x"51",
          6763 => x"82",
          6764 => x"55",
          6765 => x"51",
          6766 => x"82",
          6767 => x"83",
          6768 => x"53",
          6769 => x"80",
          6770 => x"38",
          6771 => x"78",
          6772 => x"2a",
          6773 => x"78",
          6774 => x"86",
          6775 => x"22",
          6776 => x"31",
          6777 => x"9d",
          6778 => x"98",
          6779 => x"b6",
          6780 => x"2e",
          6781 => x"82",
          6782 => x"80",
          6783 => x"f5",
          6784 => x"83",
          6785 => x"ff",
          6786 => x"38",
          6787 => x"9f",
          6788 => x"38",
          6789 => x"39",
          6790 => x"80",
          6791 => x"38",
          6792 => x"98",
          6793 => x"a0",
          6794 => x"1c",
          6795 => x"0c",
          6796 => x"17",
          6797 => x"76",
          6798 => x"81",
          6799 => x"80",
          6800 => x"d9",
          6801 => x"b6",
          6802 => x"ff",
          6803 => x"8d",
          6804 => x"8e",
          6805 => x"8a",
          6806 => x"14",
          6807 => x"3f",
          6808 => x"08",
          6809 => x"74",
          6810 => x"a2",
          6811 => x"79",
          6812 => x"ee",
          6813 => x"a8",
          6814 => x"15",
          6815 => x"2e",
          6816 => x"10",
          6817 => x"2a",
          6818 => x"05",
          6819 => x"ff",
          6820 => x"53",
          6821 => x"9c",
          6822 => x"81",
          6823 => x"0b",
          6824 => x"ff",
          6825 => x"0c",
          6826 => x"84",
          6827 => x"83",
          6828 => x"06",
          6829 => x"80",
          6830 => x"d8",
          6831 => x"b6",
          6832 => x"ff",
          6833 => x"72",
          6834 => x"81",
          6835 => x"38",
          6836 => x"73",
          6837 => x"3f",
          6838 => x"08",
          6839 => x"82",
          6840 => x"84",
          6841 => x"b2",
          6842 => x"87",
          6843 => x"98",
          6844 => x"ff",
          6845 => x"82",
          6846 => x"09",
          6847 => x"c8",
          6848 => x"51",
          6849 => x"82",
          6850 => x"84",
          6851 => x"d2",
          6852 => x"06",
          6853 => x"98",
          6854 => x"ee",
          6855 => x"98",
          6856 => x"85",
          6857 => x"09",
          6858 => x"38",
          6859 => x"51",
          6860 => x"82",
          6861 => x"90",
          6862 => x"a0",
          6863 => x"ca",
          6864 => x"98",
          6865 => x"0c",
          6866 => x"82",
          6867 => x"81",
          6868 => x"82",
          6869 => x"72",
          6870 => x"80",
          6871 => x"0c",
          6872 => x"82",
          6873 => x"90",
          6874 => x"fb",
          6875 => x"54",
          6876 => x"80",
          6877 => x"73",
          6878 => x"80",
          6879 => x"72",
          6880 => x"80",
          6881 => x"86",
          6882 => x"15",
          6883 => x"71",
          6884 => x"81",
          6885 => x"81",
          6886 => x"d0",
          6887 => x"b6",
          6888 => x"06",
          6889 => x"38",
          6890 => x"54",
          6891 => x"80",
          6892 => x"71",
          6893 => x"82",
          6894 => x"87",
          6895 => x"fa",
          6896 => x"ab",
          6897 => x"58",
          6898 => x"05",
          6899 => x"e6",
          6900 => x"80",
          6901 => x"98",
          6902 => x"38",
          6903 => x"08",
          6904 => x"cd",
          6905 => x"08",
          6906 => x"80",
          6907 => x"80",
          6908 => x"54",
          6909 => x"84",
          6910 => x"34",
          6911 => x"75",
          6912 => x"2e",
          6913 => x"53",
          6914 => x"53",
          6915 => x"f7",
          6916 => x"b6",
          6917 => x"73",
          6918 => x"0c",
          6919 => x"04",
          6920 => x"67",
          6921 => x"80",
          6922 => x"59",
          6923 => x"78",
          6924 => x"c8",
          6925 => x"06",
          6926 => x"3d",
          6927 => x"99",
          6928 => x"52",
          6929 => x"3f",
          6930 => x"08",
          6931 => x"98",
          6932 => x"38",
          6933 => x"52",
          6934 => x"52",
          6935 => x"3f",
          6936 => x"08",
          6937 => x"98",
          6938 => x"02",
          6939 => x"33",
          6940 => x"55",
          6941 => x"25",
          6942 => x"55",
          6943 => x"54",
          6944 => x"81",
          6945 => x"80",
          6946 => x"74",
          6947 => x"81",
          6948 => x"75",
          6949 => x"3f",
          6950 => x"08",
          6951 => x"02",
          6952 => x"91",
          6953 => x"81",
          6954 => x"82",
          6955 => x"06",
          6956 => x"80",
          6957 => x"88",
          6958 => x"39",
          6959 => x"58",
          6960 => x"38",
          6961 => x"70",
          6962 => x"54",
          6963 => x"81",
          6964 => x"52",
          6965 => x"a5",
          6966 => x"98",
          6967 => x"88",
          6968 => x"62",
          6969 => x"d4",
          6970 => x"54",
          6971 => x"15",
          6972 => x"62",
          6973 => x"e8",
          6974 => x"52",
          6975 => x"51",
          6976 => x"7a",
          6977 => x"83",
          6978 => x"80",
          6979 => x"38",
          6980 => x"08",
          6981 => x"53",
          6982 => x"3d",
          6983 => x"dd",
          6984 => x"b6",
          6985 => x"82",
          6986 => x"82",
          6987 => x"39",
          6988 => x"38",
          6989 => x"33",
          6990 => x"70",
          6991 => x"55",
          6992 => x"2e",
          6993 => x"55",
          6994 => x"77",
          6995 => x"81",
          6996 => x"73",
          6997 => x"38",
          6998 => x"54",
          6999 => x"a0",
          7000 => x"82",
          7001 => x"52",
          7002 => x"a3",
          7003 => x"98",
          7004 => x"18",
          7005 => x"55",
          7006 => x"98",
          7007 => x"38",
          7008 => x"70",
          7009 => x"54",
          7010 => x"86",
          7011 => x"c0",
          7012 => x"b0",
          7013 => x"1b",
          7014 => x"1b",
          7015 => x"70",
          7016 => x"d9",
          7017 => x"98",
          7018 => x"98",
          7019 => x"0c",
          7020 => x"52",
          7021 => x"3f",
          7022 => x"08",
          7023 => x"08",
          7024 => x"77",
          7025 => x"86",
          7026 => x"1a",
          7027 => x"1a",
          7028 => x"91",
          7029 => x"0b",
          7030 => x"80",
          7031 => x"0c",
          7032 => x"70",
          7033 => x"54",
          7034 => x"81",
          7035 => x"b6",
          7036 => x"2e",
          7037 => x"82",
          7038 => x"94",
          7039 => x"17",
          7040 => x"2b",
          7041 => x"57",
          7042 => x"52",
          7043 => x"9f",
          7044 => x"98",
          7045 => x"b6",
          7046 => x"26",
          7047 => x"55",
          7048 => x"08",
          7049 => x"81",
          7050 => x"79",
          7051 => x"31",
          7052 => x"70",
          7053 => x"25",
          7054 => x"76",
          7055 => x"81",
          7056 => x"55",
          7057 => x"38",
          7058 => x"0c",
          7059 => x"75",
          7060 => x"54",
          7061 => x"a2",
          7062 => x"7a",
          7063 => x"3f",
          7064 => x"08",
          7065 => x"55",
          7066 => x"89",
          7067 => x"98",
          7068 => x"1a",
          7069 => x"80",
          7070 => x"54",
          7071 => x"98",
          7072 => x"0d",
          7073 => x"0d",
          7074 => x"64",
          7075 => x"59",
          7076 => x"90",
          7077 => x"52",
          7078 => x"cf",
          7079 => x"98",
          7080 => x"b6",
          7081 => x"38",
          7082 => x"55",
          7083 => x"86",
          7084 => x"82",
          7085 => x"19",
          7086 => x"55",
          7087 => x"80",
          7088 => x"38",
          7089 => x"0b",
          7090 => x"82",
          7091 => x"39",
          7092 => x"1a",
          7093 => x"82",
          7094 => x"19",
          7095 => x"08",
          7096 => x"7c",
          7097 => x"74",
          7098 => x"2e",
          7099 => x"94",
          7100 => x"83",
          7101 => x"56",
          7102 => x"38",
          7103 => x"22",
          7104 => x"89",
          7105 => x"55",
          7106 => x"75",
          7107 => x"19",
          7108 => x"39",
          7109 => x"52",
          7110 => x"93",
          7111 => x"98",
          7112 => x"75",
          7113 => x"38",
          7114 => x"ff",
          7115 => x"98",
          7116 => x"19",
          7117 => x"51",
          7118 => x"82",
          7119 => x"80",
          7120 => x"38",
          7121 => x"08",
          7122 => x"2a",
          7123 => x"80",
          7124 => x"38",
          7125 => x"8a",
          7126 => x"5c",
          7127 => x"27",
          7128 => x"7a",
          7129 => x"54",
          7130 => x"52",
          7131 => x"51",
          7132 => x"82",
          7133 => x"fe",
          7134 => x"83",
          7135 => x"56",
          7136 => x"9f",
          7137 => x"08",
          7138 => x"74",
          7139 => x"38",
          7140 => x"b4",
          7141 => x"16",
          7142 => x"89",
          7143 => x"51",
          7144 => x"77",
          7145 => x"b9",
          7146 => x"1a",
          7147 => x"08",
          7148 => x"84",
          7149 => x"57",
          7150 => x"27",
          7151 => x"56",
          7152 => x"52",
          7153 => x"c7",
          7154 => x"98",
          7155 => x"38",
          7156 => x"19",
          7157 => x"06",
          7158 => x"52",
          7159 => x"a2",
          7160 => x"31",
          7161 => x"7f",
          7162 => x"94",
          7163 => x"94",
          7164 => x"5c",
          7165 => x"80",
          7166 => x"b6",
          7167 => x"3d",
          7168 => x"3d",
          7169 => x"65",
          7170 => x"5d",
          7171 => x"0c",
          7172 => x"05",
          7173 => x"f6",
          7174 => x"b6",
          7175 => x"82",
          7176 => x"8a",
          7177 => x"33",
          7178 => x"2e",
          7179 => x"56",
          7180 => x"90",
          7181 => x"81",
          7182 => x"06",
          7183 => x"87",
          7184 => x"2e",
          7185 => x"95",
          7186 => x"91",
          7187 => x"56",
          7188 => x"81",
          7189 => x"34",
          7190 => x"8e",
          7191 => x"08",
          7192 => x"56",
          7193 => x"84",
          7194 => x"5c",
          7195 => x"82",
          7196 => x"18",
          7197 => x"ff",
          7198 => x"74",
          7199 => x"7e",
          7200 => x"ff",
          7201 => x"2a",
          7202 => x"7a",
          7203 => x"8c",
          7204 => x"08",
          7205 => x"38",
          7206 => x"39",
          7207 => x"52",
          7208 => x"e7",
          7209 => x"98",
          7210 => x"b6",
          7211 => x"2e",
          7212 => x"74",
          7213 => x"91",
          7214 => x"2e",
          7215 => x"74",
          7216 => x"88",
          7217 => x"38",
          7218 => x"0c",
          7219 => x"15",
          7220 => x"08",
          7221 => x"06",
          7222 => x"51",
          7223 => x"82",
          7224 => x"fe",
          7225 => x"18",
          7226 => x"51",
          7227 => x"82",
          7228 => x"80",
          7229 => x"38",
          7230 => x"08",
          7231 => x"2a",
          7232 => x"80",
          7233 => x"38",
          7234 => x"8a",
          7235 => x"5b",
          7236 => x"27",
          7237 => x"7b",
          7238 => x"54",
          7239 => x"52",
          7240 => x"51",
          7241 => x"82",
          7242 => x"fe",
          7243 => x"b0",
          7244 => x"31",
          7245 => x"79",
          7246 => x"84",
          7247 => x"16",
          7248 => x"89",
          7249 => x"52",
          7250 => x"cc",
          7251 => x"55",
          7252 => x"16",
          7253 => x"2b",
          7254 => x"39",
          7255 => x"94",
          7256 => x"93",
          7257 => x"cd",
          7258 => x"b6",
          7259 => x"e3",
          7260 => x"b0",
          7261 => x"76",
          7262 => x"94",
          7263 => x"ff",
          7264 => x"71",
          7265 => x"7b",
          7266 => x"38",
          7267 => x"18",
          7268 => x"51",
          7269 => x"82",
          7270 => x"fd",
          7271 => x"53",
          7272 => x"18",
          7273 => x"06",
          7274 => x"51",
          7275 => x"7e",
          7276 => x"83",
          7277 => x"76",
          7278 => x"17",
          7279 => x"1e",
          7280 => x"18",
          7281 => x"0c",
          7282 => x"58",
          7283 => x"74",
          7284 => x"38",
          7285 => x"8c",
          7286 => x"90",
          7287 => x"33",
          7288 => x"55",
          7289 => x"34",
          7290 => x"82",
          7291 => x"90",
          7292 => x"f8",
          7293 => x"8b",
          7294 => x"53",
          7295 => x"f2",
          7296 => x"b6",
          7297 => x"82",
          7298 => x"80",
          7299 => x"16",
          7300 => x"2a",
          7301 => x"51",
          7302 => x"80",
          7303 => x"38",
          7304 => x"52",
          7305 => x"e7",
          7306 => x"98",
          7307 => x"b6",
          7308 => x"d4",
          7309 => x"08",
          7310 => x"a0",
          7311 => x"73",
          7312 => x"88",
          7313 => x"74",
          7314 => x"51",
          7315 => x"8c",
          7316 => x"9c",
          7317 => x"fb",
          7318 => x"b2",
          7319 => x"15",
          7320 => x"3f",
          7321 => x"15",
          7322 => x"3f",
          7323 => x"0b",
          7324 => x"78",
          7325 => x"3f",
          7326 => x"08",
          7327 => x"81",
          7328 => x"57",
          7329 => x"34",
          7330 => x"98",
          7331 => x"0d",
          7332 => x"0d",
          7333 => x"54",
          7334 => x"82",
          7335 => x"53",
          7336 => x"08",
          7337 => x"3d",
          7338 => x"73",
          7339 => x"3f",
          7340 => x"08",
          7341 => x"98",
          7342 => x"82",
          7343 => x"74",
          7344 => x"b6",
          7345 => x"3d",
          7346 => x"3d",
          7347 => x"51",
          7348 => x"8b",
          7349 => x"82",
          7350 => x"24",
          7351 => x"b6",
          7352 => x"cd",
          7353 => x"52",
          7354 => x"98",
          7355 => x"0d",
          7356 => x"0d",
          7357 => x"3d",
          7358 => x"94",
          7359 => x"c1",
          7360 => x"98",
          7361 => x"b6",
          7362 => x"e0",
          7363 => x"63",
          7364 => x"d4",
          7365 => x"8d",
          7366 => x"98",
          7367 => x"b6",
          7368 => x"38",
          7369 => x"05",
          7370 => x"2b",
          7371 => x"80",
          7372 => x"76",
          7373 => x"0c",
          7374 => x"02",
          7375 => x"70",
          7376 => x"81",
          7377 => x"56",
          7378 => x"9e",
          7379 => x"53",
          7380 => x"db",
          7381 => x"b6",
          7382 => x"15",
          7383 => x"82",
          7384 => x"84",
          7385 => x"06",
          7386 => x"55",
          7387 => x"98",
          7388 => x"0d",
          7389 => x"0d",
          7390 => x"5b",
          7391 => x"80",
          7392 => x"ff",
          7393 => x"9f",
          7394 => x"b5",
          7395 => x"98",
          7396 => x"b6",
          7397 => x"fc",
          7398 => x"7a",
          7399 => x"08",
          7400 => x"64",
          7401 => x"2e",
          7402 => x"a0",
          7403 => x"70",
          7404 => x"ea",
          7405 => x"98",
          7406 => x"b6",
          7407 => x"d4",
          7408 => x"7b",
          7409 => x"3f",
          7410 => x"08",
          7411 => x"98",
          7412 => x"38",
          7413 => x"51",
          7414 => x"82",
          7415 => x"45",
          7416 => x"51",
          7417 => x"82",
          7418 => x"57",
          7419 => x"08",
          7420 => x"80",
          7421 => x"da",
          7422 => x"b6",
          7423 => x"82",
          7424 => x"a4",
          7425 => x"7b",
          7426 => x"3f",
          7427 => x"98",
          7428 => x"38",
          7429 => x"51",
          7430 => x"82",
          7431 => x"57",
          7432 => x"08",
          7433 => x"38",
          7434 => x"09",
          7435 => x"38",
          7436 => x"e0",
          7437 => x"dc",
          7438 => x"ff",
          7439 => x"74",
          7440 => x"3f",
          7441 => x"78",
          7442 => x"33",
          7443 => x"56",
          7444 => x"91",
          7445 => x"05",
          7446 => x"81",
          7447 => x"56",
          7448 => x"f5",
          7449 => x"54",
          7450 => x"81",
          7451 => x"80",
          7452 => x"78",
          7453 => x"55",
          7454 => x"11",
          7455 => x"18",
          7456 => x"58",
          7457 => x"34",
          7458 => x"ff",
          7459 => x"55",
          7460 => x"34",
          7461 => x"77",
          7462 => x"81",
          7463 => x"ff",
          7464 => x"55",
          7465 => x"34",
          7466 => x"cd",
          7467 => x"84",
          7468 => x"d0",
          7469 => x"70",
          7470 => x"56",
          7471 => x"76",
          7472 => x"81",
          7473 => x"70",
          7474 => x"56",
          7475 => x"82",
          7476 => x"78",
          7477 => x"80",
          7478 => x"27",
          7479 => x"19",
          7480 => x"7a",
          7481 => x"5c",
          7482 => x"55",
          7483 => x"7a",
          7484 => x"5c",
          7485 => x"2e",
          7486 => x"85",
          7487 => x"94",
          7488 => x"81",
          7489 => x"73",
          7490 => x"81",
          7491 => x"7a",
          7492 => x"38",
          7493 => x"76",
          7494 => x"0c",
          7495 => x"04",
          7496 => x"7b",
          7497 => x"fc",
          7498 => x"53",
          7499 => x"bb",
          7500 => x"98",
          7501 => x"b6",
          7502 => x"fa",
          7503 => x"33",
          7504 => x"f2",
          7505 => x"08",
          7506 => x"27",
          7507 => x"15",
          7508 => x"2a",
          7509 => x"51",
          7510 => x"83",
          7511 => x"94",
          7512 => x"80",
          7513 => x"0c",
          7514 => x"2e",
          7515 => x"79",
          7516 => x"70",
          7517 => x"51",
          7518 => x"2e",
          7519 => x"52",
          7520 => x"fe",
          7521 => x"82",
          7522 => x"ff",
          7523 => x"70",
          7524 => x"fe",
          7525 => x"82",
          7526 => x"73",
          7527 => x"76",
          7528 => x"06",
          7529 => x"0c",
          7530 => x"98",
          7531 => x"58",
          7532 => x"39",
          7533 => x"54",
          7534 => x"73",
          7535 => x"cd",
          7536 => x"b6",
          7537 => x"82",
          7538 => x"81",
          7539 => x"38",
          7540 => x"08",
          7541 => x"9b",
          7542 => x"98",
          7543 => x"0c",
          7544 => x"0c",
          7545 => x"81",
          7546 => x"76",
          7547 => x"38",
          7548 => x"94",
          7549 => x"94",
          7550 => x"16",
          7551 => x"2a",
          7552 => x"51",
          7553 => x"72",
          7554 => x"38",
          7555 => x"51",
          7556 => x"82",
          7557 => x"54",
          7558 => x"08",
          7559 => x"b6",
          7560 => x"a7",
          7561 => x"74",
          7562 => x"3f",
          7563 => x"08",
          7564 => x"2e",
          7565 => x"74",
          7566 => x"79",
          7567 => x"14",
          7568 => x"38",
          7569 => x"0c",
          7570 => x"94",
          7571 => x"94",
          7572 => x"83",
          7573 => x"72",
          7574 => x"38",
          7575 => x"51",
          7576 => x"82",
          7577 => x"94",
          7578 => x"91",
          7579 => x"53",
          7580 => x"81",
          7581 => x"34",
          7582 => x"39",
          7583 => x"82",
          7584 => x"05",
          7585 => x"08",
          7586 => x"08",
          7587 => x"38",
          7588 => x"0c",
          7589 => x"80",
          7590 => x"72",
          7591 => x"73",
          7592 => x"53",
          7593 => x"8c",
          7594 => x"16",
          7595 => x"38",
          7596 => x"0c",
          7597 => x"82",
          7598 => x"8b",
          7599 => x"f9",
          7600 => x"56",
          7601 => x"80",
          7602 => x"38",
          7603 => x"3d",
          7604 => x"8a",
          7605 => x"51",
          7606 => x"82",
          7607 => x"55",
          7608 => x"08",
          7609 => x"77",
          7610 => x"52",
          7611 => x"b5",
          7612 => x"98",
          7613 => x"b6",
          7614 => x"c3",
          7615 => x"33",
          7616 => x"55",
          7617 => x"24",
          7618 => x"16",
          7619 => x"2a",
          7620 => x"51",
          7621 => x"80",
          7622 => x"9c",
          7623 => x"77",
          7624 => x"3f",
          7625 => x"08",
          7626 => x"77",
          7627 => x"22",
          7628 => x"74",
          7629 => x"ce",
          7630 => x"b6",
          7631 => x"74",
          7632 => x"81",
          7633 => x"85",
          7634 => x"74",
          7635 => x"38",
          7636 => x"74",
          7637 => x"b6",
          7638 => x"3d",
          7639 => x"3d",
          7640 => x"3d",
          7641 => x"70",
          7642 => x"ff",
          7643 => x"98",
          7644 => x"82",
          7645 => x"73",
          7646 => x"0d",
          7647 => x"0d",
          7648 => x"3d",
          7649 => x"71",
          7650 => x"e7",
          7651 => x"b6",
          7652 => x"82",
          7653 => x"80",
          7654 => x"93",
          7655 => x"98",
          7656 => x"51",
          7657 => x"82",
          7658 => x"53",
          7659 => x"82",
          7660 => x"52",
          7661 => x"ac",
          7662 => x"98",
          7663 => x"b6",
          7664 => x"2e",
          7665 => x"85",
          7666 => x"87",
          7667 => x"98",
          7668 => x"74",
          7669 => x"d5",
          7670 => x"52",
          7671 => x"89",
          7672 => x"98",
          7673 => x"70",
          7674 => x"07",
          7675 => x"82",
          7676 => x"06",
          7677 => x"54",
          7678 => x"98",
          7679 => x"0d",
          7680 => x"0d",
          7681 => x"53",
          7682 => x"53",
          7683 => x"56",
          7684 => x"82",
          7685 => x"55",
          7686 => x"08",
          7687 => x"52",
          7688 => x"81",
          7689 => x"98",
          7690 => x"b6",
          7691 => x"38",
          7692 => x"05",
          7693 => x"2b",
          7694 => x"80",
          7695 => x"86",
          7696 => x"76",
          7697 => x"38",
          7698 => x"51",
          7699 => x"74",
          7700 => x"0c",
          7701 => x"04",
          7702 => x"63",
          7703 => x"80",
          7704 => x"ec",
          7705 => x"3d",
          7706 => x"3f",
          7707 => x"08",
          7708 => x"98",
          7709 => x"38",
          7710 => x"73",
          7711 => x"08",
          7712 => x"13",
          7713 => x"58",
          7714 => x"26",
          7715 => x"7c",
          7716 => x"39",
          7717 => x"cc",
          7718 => x"81",
          7719 => x"b6",
          7720 => x"33",
          7721 => x"81",
          7722 => x"06",
          7723 => x"75",
          7724 => x"52",
          7725 => x"05",
          7726 => x"3f",
          7727 => x"08",
          7728 => x"38",
          7729 => x"08",
          7730 => x"38",
          7731 => x"08",
          7732 => x"b6",
          7733 => x"80",
          7734 => x"81",
          7735 => x"59",
          7736 => x"14",
          7737 => x"ca",
          7738 => x"39",
          7739 => x"82",
          7740 => x"57",
          7741 => x"38",
          7742 => x"18",
          7743 => x"ff",
          7744 => x"82",
          7745 => x"5b",
          7746 => x"08",
          7747 => x"7c",
          7748 => x"12",
          7749 => x"52",
          7750 => x"82",
          7751 => x"06",
          7752 => x"14",
          7753 => x"cb",
          7754 => x"98",
          7755 => x"ff",
          7756 => x"70",
          7757 => x"82",
          7758 => x"51",
          7759 => x"b4",
          7760 => x"bb",
          7761 => x"b6",
          7762 => x"0a",
          7763 => x"70",
          7764 => x"84",
          7765 => x"51",
          7766 => x"ff",
          7767 => x"56",
          7768 => x"38",
          7769 => x"7c",
          7770 => x"0c",
          7771 => x"81",
          7772 => x"74",
          7773 => x"7a",
          7774 => x"0c",
          7775 => x"04",
          7776 => x"79",
          7777 => x"05",
          7778 => x"57",
          7779 => x"82",
          7780 => x"56",
          7781 => x"08",
          7782 => x"91",
          7783 => x"75",
          7784 => x"90",
          7785 => x"81",
          7786 => x"06",
          7787 => x"87",
          7788 => x"2e",
          7789 => x"94",
          7790 => x"73",
          7791 => x"27",
          7792 => x"73",
          7793 => x"b6",
          7794 => x"88",
          7795 => x"76",
          7796 => x"3f",
          7797 => x"08",
          7798 => x"0c",
          7799 => x"39",
          7800 => x"52",
          7801 => x"bf",
          7802 => x"b6",
          7803 => x"2e",
          7804 => x"83",
          7805 => x"82",
          7806 => x"81",
          7807 => x"06",
          7808 => x"56",
          7809 => x"a0",
          7810 => x"82",
          7811 => x"98",
          7812 => x"94",
          7813 => x"08",
          7814 => x"98",
          7815 => x"51",
          7816 => x"82",
          7817 => x"56",
          7818 => x"8c",
          7819 => x"17",
          7820 => x"07",
          7821 => x"18",
          7822 => x"2e",
          7823 => x"91",
          7824 => x"55",
          7825 => x"98",
          7826 => x"0d",
          7827 => x"0d",
          7828 => x"3d",
          7829 => x"52",
          7830 => x"da",
          7831 => x"b6",
          7832 => x"82",
          7833 => x"81",
          7834 => x"45",
          7835 => x"52",
          7836 => x"52",
          7837 => x"3f",
          7838 => x"08",
          7839 => x"98",
          7840 => x"38",
          7841 => x"05",
          7842 => x"2a",
          7843 => x"51",
          7844 => x"55",
          7845 => x"38",
          7846 => x"54",
          7847 => x"81",
          7848 => x"80",
          7849 => x"70",
          7850 => x"54",
          7851 => x"81",
          7852 => x"52",
          7853 => x"c5",
          7854 => x"98",
          7855 => x"2a",
          7856 => x"51",
          7857 => x"80",
          7858 => x"38",
          7859 => x"b6",
          7860 => x"15",
          7861 => x"86",
          7862 => x"82",
          7863 => x"5c",
          7864 => x"3d",
          7865 => x"c7",
          7866 => x"b6",
          7867 => x"82",
          7868 => x"80",
          7869 => x"b6",
          7870 => x"73",
          7871 => x"3f",
          7872 => x"08",
          7873 => x"98",
          7874 => x"87",
          7875 => x"39",
          7876 => x"08",
          7877 => x"38",
          7878 => x"08",
          7879 => x"77",
          7880 => x"3f",
          7881 => x"08",
          7882 => x"08",
          7883 => x"b6",
          7884 => x"80",
          7885 => x"55",
          7886 => x"94",
          7887 => x"2e",
          7888 => x"53",
          7889 => x"51",
          7890 => x"82",
          7891 => x"55",
          7892 => x"78",
          7893 => x"fe",
          7894 => x"98",
          7895 => x"82",
          7896 => x"a0",
          7897 => x"e9",
          7898 => x"53",
          7899 => x"05",
          7900 => x"51",
          7901 => x"82",
          7902 => x"54",
          7903 => x"08",
          7904 => x"78",
          7905 => x"8e",
          7906 => x"58",
          7907 => x"82",
          7908 => x"54",
          7909 => x"08",
          7910 => x"54",
          7911 => x"82",
          7912 => x"84",
          7913 => x"06",
          7914 => x"02",
          7915 => x"33",
          7916 => x"81",
          7917 => x"86",
          7918 => x"f6",
          7919 => x"74",
          7920 => x"70",
          7921 => x"c3",
          7922 => x"98",
          7923 => x"56",
          7924 => x"08",
          7925 => x"54",
          7926 => x"08",
          7927 => x"81",
          7928 => x"82",
          7929 => x"98",
          7930 => x"09",
          7931 => x"38",
          7932 => x"b4",
          7933 => x"b0",
          7934 => x"98",
          7935 => x"51",
          7936 => x"82",
          7937 => x"54",
          7938 => x"08",
          7939 => x"8b",
          7940 => x"b4",
          7941 => x"b7",
          7942 => x"54",
          7943 => x"15",
          7944 => x"90",
          7945 => x"34",
          7946 => x"0a",
          7947 => x"19",
          7948 => x"9f",
          7949 => x"78",
          7950 => x"51",
          7951 => x"a0",
          7952 => x"11",
          7953 => x"05",
          7954 => x"b6",
          7955 => x"ae",
          7956 => x"15",
          7957 => x"78",
          7958 => x"53",
          7959 => x"3f",
          7960 => x"0b",
          7961 => x"77",
          7962 => x"3f",
          7963 => x"08",
          7964 => x"98",
          7965 => x"82",
          7966 => x"52",
          7967 => x"51",
          7968 => x"3f",
          7969 => x"52",
          7970 => x"aa",
          7971 => x"90",
          7972 => x"34",
          7973 => x"0b",
          7974 => x"78",
          7975 => x"b6",
          7976 => x"98",
          7977 => x"39",
          7978 => x"52",
          7979 => x"be",
          7980 => x"82",
          7981 => x"99",
          7982 => x"da",
          7983 => x"3d",
          7984 => x"d2",
          7985 => x"53",
          7986 => x"84",
          7987 => x"3d",
          7988 => x"3f",
          7989 => x"08",
          7990 => x"98",
          7991 => x"38",
          7992 => x"3d",
          7993 => x"3d",
          7994 => x"cc",
          7995 => x"b6",
          7996 => x"82",
          7997 => x"82",
          7998 => x"81",
          7999 => x"81",
          8000 => x"86",
          8001 => x"aa",
          8002 => x"a4",
          8003 => x"a8",
          8004 => x"05",
          8005 => x"ea",
          8006 => x"77",
          8007 => x"70",
          8008 => x"b4",
          8009 => x"3d",
          8010 => x"51",
          8011 => x"82",
          8012 => x"55",
          8013 => x"08",
          8014 => x"6f",
          8015 => x"06",
          8016 => x"a2",
          8017 => x"92",
          8018 => x"81",
          8019 => x"b6",
          8020 => x"2e",
          8021 => x"81",
          8022 => x"51",
          8023 => x"82",
          8024 => x"55",
          8025 => x"08",
          8026 => x"68",
          8027 => x"a8",
          8028 => x"05",
          8029 => x"51",
          8030 => x"3f",
          8031 => x"33",
          8032 => x"8b",
          8033 => x"84",
          8034 => x"06",
          8035 => x"73",
          8036 => x"a0",
          8037 => x"8b",
          8038 => x"54",
          8039 => x"15",
          8040 => x"33",
          8041 => x"70",
          8042 => x"55",
          8043 => x"2e",
          8044 => x"6e",
          8045 => x"df",
          8046 => x"78",
          8047 => x"3f",
          8048 => x"08",
          8049 => x"ff",
          8050 => x"82",
          8051 => x"98",
          8052 => x"80",
          8053 => x"b6",
          8054 => x"78",
          8055 => x"af",
          8056 => x"98",
          8057 => x"d4",
          8058 => x"55",
          8059 => x"08",
          8060 => x"81",
          8061 => x"73",
          8062 => x"81",
          8063 => x"63",
          8064 => x"76",
          8065 => x"3f",
          8066 => x"0b",
          8067 => x"87",
          8068 => x"98",
          8069 => x"77",
          8070 => x"3f",
          8071 => x"08",
          8072 => x"98",
          8073 => x"78",
          8074 => x"aa",
          8075 => x"98",
          8076 => x"82",
          8077 => x"a8",
          8078 => x"ed",
          8079 => x"80",
          8080 => x"02",
          8081 => x"df",
          8082 => x"57",
          8083 => x"3d",
          8084 => x"96",
          8085 => x"e9",
          8086 => x"98",
          8087 => x"b6",
          8088 => x"cf",
          8089 => x"65",
          8090 => x"d4",
          8091 => x"b5",
          8092 => x"98",
          8093 => x"b6",
          8094 => x"38",
          8095 => x"05",
          8096 => x"06",
          8097 => x"73",
          8098 => x"a7",
          8099 => x"09",
          8100 => x"71",
          8101 => x"06",
          8102 => x"55",
          8103 => x"15",
          8104 => x"81",
          8105 => x"34",
          8106 => x"b4",
          8107 => x"b6",
          8108 => x"74",
          8109 => x"0c",
          8110 => x"04",
          8111 => x"64",
          8112 => x"93",
          8113 => x"52",
          8114 => x"d1",
          8115 => x"b6",
          8116 => x"82",
          8117 => x"80",
          8118 => x"58",
          8119 => x"3d",
          8120 => x"c8",
          8121 => x"b6",
          8122 => x"82",
          8123 => x"b4",
          8124 => x"c7",
          8125 => x"a0",
          8126 => x"55",
          8127 => x"84",
          8128 => x"17",
          8129 => x"2b",
          8130 => x"96",
          8131 => x"b0",
          8132 => x"54",
          8133 => x"15",
          8134 => x"ff",
          8135 => x"82",
          8136 => x"55",
          8137 => x"98",
          8138 => x"0d",
          8139 => x"0d",
          8140 => x"5a",
          8141 => x"3d",
          8142 => x"99",
          8143 => x"81",
          8144 => x"98",
          8145 => x"98",
          8146 => x"82",
          8147 => x"07",
          8148 => x"55",
          8149 => x"2e",
          8150 => x"81",
          8151 => x"55",
          8152 => x"2e",
          8153 => x"7b",
          8154 => x"80",
          8155 => x"70",
          8156 => x"be",
          8157 => x"b6",
          8158 => x"82",
          8159 => x"80",
          8160 => x"52",
          8161 => x"dc",
          8162 => x"98",
          8163 => x"b6",
          8164 => x"38",
          8165 => x"08",
          8166 => x"08",
          8167 => x"56",
          8168 => x"19",
          8169 => x"59",
          8170 => x"74",
          8171 => x"56",
          8172 => x"ec",
          8173 => x"75",
          8174 => x"74",
          8175 => x"2e",
          8176 => x"16",
          8177 => x"33",
          8178 => x"73",
          8179 => x"38",
          8180 => x"84",
          8181 => x"06",
          8182 => x"7a",
          8183 => x"76",
          8184 => x"07",
          8185 => x"54",
          8186 => x"80",
          8187 => x"80",
          8188 => x"7b",
          8189 => x"53",
          8190 => x"93",
          8191 => x"98",
          8192 => x"b6",
          8193 => x"38",
          8194 => x"55",
          8195 => x"56",
          8196 => x"8b",
          8197 => x"56",
          8198 => x"83",
          8199 => x"75",
          8200 => x"51",
          8201 => x"3f",
          8202 => x"08",
          8203 => x"82",
          8204 => x"98",
          8205 => x"e6",
          8206 => x"53",
          8207 => x"b8",
          8208 => x"3d",
          8209 => x"3f",
          8210 => x"08",
          8211 => x"08",
          8212 => x"b6",
          8213 => x"98",
          8214 => x"a0",
          8215 => x"70",
          8216 => x"ae",
          8217 => x"6d",
          8218 => x"81",
          8219 => x"57",
          8220 => x"74",
          8221 => x"38",
          8222 => x"81",
          8223 => x"81",
          8224 => x"52",
          8225 => x"89",
          8226 => x"98",
          8227 => x"a5",
          8228 => x"33",
          8229 => x"54",
          8230 => x"3f",
          8231 => x"08",
          8232 => x"38",
          8233 => x"76",
          8234 => x"05",
          8235 => x"39",
          8236 => x"08",
          8237 => x"15",
          8238 => x"ff",
          8239 => x"73",
          8240 => x"38",
          8241 => x"83",
          8242 => x"56",
          8243 => x"75",
          8244 => x"82",
          8245 => x"33",
          8246 => x"2e",
          8247 => x"52",
          8248 => x"51",
          8249 => x"3f",
          8250 => x"08",
          8251 => x"ff",
          8252 => x"38",
          8253 => x"88",
          8254 => x"8a",
          8255 => x"38",
          8256 => x"ec",
          8257 => x"75",
          8258 => x"74",
          8259 => x"73",
          8260 => x"05",
          8261 => x"17",
          8262 => x"70",
          8263 => x"34",
          8264 => x"70",
          8265 => x"ff",
          8266 => x"55",
          8267 => x"26",
          8268 => x"8b",
          8269 => x"86",
          8270 => x"e5",
          8271 => x"38",
          8272 => x"99",
          8273 => x"05",
          8274 => x"70",
          8275 => x"73",
          8276 => x"81",
          8277 => x"ff",
          8278 => x"ed",
          8279 => x"80",
          8280 => x"91",
          8281 => x"55",
          8282 => x"3f",
          8283 => x"08",
          8284 => x"98",
          8285 => x"38",
          8286 => x"51",
          8287 => x"3f",
          8288 => x"08",
          8289 => x"98",
          8290 => x"76",
          8291 => x"67",
          8292 => x"34",
          8293 => x"82",
          8294 => x"84",
          8295 => x"06",
          8296 => x"80",
          8297 => x"2e",
          8298 => x"81",
          8299 => x"ff",
          8300 => x"82",
          8301 => x"54",
          8302 => x"08",
          8303 => x"53",
          8304 => x"08",
          8305 => x"ff",
          8306 => x"67",
          8307 => x"8b",
          8308 => x"53",
          8309 => x"51",
          8310 => x"3f",
          8311 => x"0b",
          8312 => x"79",
          8313 => x"ee",
          8314 => x"98",
          8315 => x"55",
          8316 => x"98",
          8317 => x"0d",
          8318 => x"0d",
          8319 => x"88",
          8320 => x"05",
          8321 => x"fc",
          8322 => x"54",
          8323 => x"d2",
          8324 => x"b6",
          8325 => x"82",
          8326 => x"82",
          8327 => x"1a",
          8328 => x"82",
          8329 => x"80",
          8330 => x"8c",
          8331 => x"78",
          8332 => x"1a",
          8333 => x"2a",
          8334 => x"51",
          8335 => x"90",
          8336 => x"82",
          8337 => x"58",
          8338 => x"81",
          8339 => x"39",
          8340 => x"22",
          8341 => x"70",
          8342 => x"56",
          8343 => x"c2",
          8344 => x"14",
          8345 => x"30",
          8346 => x"9f",
          8347 => x"98",
          8348 => x"19",
          8349 => x"5a",
          8350 => x"81",
          8351 => x"38",
          8352 => x"77",
          8353 => x"82",
          8354 => x"56",
          8355 => x"74",
          8356 => x"ff",
          8357 => x"81",
          8358 => x"55",
          8359 => x"75",
          8360 => x"82",
          8361 => x"98",
          8362 => x"ff",
          8363 => x"b6",
          8364 => x"2e",
          8365 => x"82",
          8366 => x"8e",
          8367 => x"56",
          8368 => x"09",
          8369 => x"38",
          8370 => x"59",
          8371 => x"77",
          8372 => x"06",
          8373 => x"87",
          8374 => x"39",
          8375 => x"ba",
          8376 => x"55",
          8377 => x"2e",
          8378 => x"15",
          8379 => x"2e",
          8380 => x"83",
          8381 => x"75",
          8382 => x"7e",
          8383 => x"a8",
          8384 => x"98",
          8385 => x"b6",
          8386 => x"ce",
          8387 => x"16",
          8388 => x"56",
          8389 => x"38",
          8390 => x"19",
          8391 => x"8c",
          8392 => x"7d",
          8393 => x"38",
          8394 => x"0c",
          8395 => x"0c",
          8396 => x"80",
          8397 => x"73",
          8398 => x"98",
          8399 => x"05",
          8400 => x"57",
          8401 => x"26",
          8402 => x"7b",
          8403 => x"0c",
          8404 => x"81",
          8405 => x"84",
          8406 => x"54",
          8407 => x"98",
          8408 => x"0d",
          8409 => x"0d",
          8410 => x"88",
          8411 => x"05",
          8412 => x"54",
          8413 => x"c5",
          8414 => x"56",
          8415 => x"b6",
          8416 => x"8b",
          8417 => x"b6",
          8418 => x"29",
          8419 => x"05",
          8420 => x"55",
          8421 => x"84",
          8422 => x"34",
          8423 => x"08",
          8424 => x"5f",
          8425 => x"51",
          8426 => x"3f",
          8427 => x"08",
          8428 => x"70",
          8429 => x"57",
          8430 => x"8b",
          8431 => x"82",
          8432 => x"06",
          8433 => x"56",
          8434 => x"38",
          8435 => x"05",
          8436 => x"7e",
          8437 => x"f0",
          8438 => x"98",
          8439 => x"67",
          8440 => x"2e",
          8441 => x"82",
          8442 => x"8b",
          8443 => x"75",
          8444 => x"80",
          8445 => x"81",
          8446 => x"2e",
          8447 => x"80",
          8448 => x"38",
          8449 => x"0a",
          8450 => x"ff",
          8451 => x"55",
          8452 => x"86",
          8453 => x"8a",
          8454 => x"89",
          8455 => x"2a",
          8456 => x"77",
          8457 => x"59",
          8458 => x"81",
          8459 => x"70",
          8460 => x"07",
          8461 => x"56",
          8462 => x"38",
          8463 => x"05",
          8464 => x"7e",
          8465 => x"80",
          8466 => x"82",
          8467 => x"8a",
          8468 => x"83",
          8469 => x"06",
          8470 => x"08",
          8471 => x"74",
          8472 => x"41",
          8473 => x"56",
          8474 => x"8a",
          8475 => x"61",
          8476 => x"55",
          8477 => x"27",
          8478 => x"93",
          8479 => x"80",
          8480 => x"38",
          8481 => x"70",
          8482 => x"43",
          8483 => x"95",
          8484 => x"06",
          8485 => x"2e",
          8486 => x"77",
          8487 => x"74",
          8488 => x"83",
          8489 => x"06",
          8490 => x"82",
          8491 => x"2e",
          8492 => x"78",
          8493 => x"2e",
          8494 => x"80",
          8495 => x"ae",
          8496 => x"2a",
          8497 => x"82",
          8498 => x"56",
          8499 => x"2e",
          8500 => x"77",
          8501 => x"82",
          8502 => x"79",
          8503 => x"70",
          8504 => x"5a",
          8505 => x"86",
          8506 => x"27",
          8507 => x"52",
          8508 => x"bd",
          8509 => x"b6",
          8510 => x"29",
          8511 => x"70",
          8512 => x"55",
          8513 => x"0b",
          8514 => x"08",
          8515 => x"05",
          8516 => x"ff",
          8517 => x"27",
          8518 => x"88",
          8519 => x"ae",
          8520 => x"2a",
          8521 => x"82",
          8522 => x"56",
          8523 => x"2e",
          8524 => x"77",
          8525 => x"82",
          8526 => x"79",
          8527 => x"70",
          8528 => x"5a",
          8529 => x"86",
          8530 => x"27",
          8531 => x"52",
          8532 => x"bc",
          8533 => x"b6",
          8534 => x"84",
          8535 => x"b6",
          8536 => x"f5",
          8537 => x"81",
          8538 => x"98",
          8539 => x"b6",
          8540 => x"71",
          8541 => x"83",
          8542 => x"5e",
          8543 => x"89",
          8544 => x"5c",
          8545 => x"1c",
          8546 => x"05",
          8547 => x"ff",
          8548 => x"70",
          8549 => x"31",
          8550 => x"57",
          8551 => x"83",
          8552 => x"06",
          8553 => x"1c",
          8554 => x"5c",
          8555 => x"1d",
          8556 => x"29",
          8557 => x"31",
          8558 => x"55",
          8559 => x"87",
          8560 => x"7c",
          8561 => x"7a",
          8562 => x"31",
          8563 => x"bb",
          8564 => x"b6",
          8565 => x"7d",
          8566 => x"81",
          8567 => x"82",
          8568 => x"83",
          8569 => x"80",
          8570 => x"87",
          8571 => x"81",
          8572 => x"fd",
          8573 => x"f8",
          8574 => x"2e",
          8575 => x"80",
          8576 => x"ff",
          8577 => x"b6",
          8578 => x"a0",
          8579 => x"38",
          8580 => x"74",
          8581 => x"86",
          8582 => x"fd",
          8583 => x"81",
          8584 => x"80",
          8585 => x"83",
          8586 => x"39",
          8587 => x"08",
          8588 => x"92",
          8589 => x"b8",
          8590 => x"59",
          8591 => x"27",
          8592 => x"86",
          8593 => x"55",
          8594 => x"09",
          8595 => x"38",
          8596 => x"f5",
          8597 => x"38",
          8598 => x"55",
          8599 => x"86",
          8600 => x"80",
          8601 => x"7a",
          8602 => x"b9",
          8603 => x"82",
          8604 => x"7a",
          8605 => x"8a",
          8606 => x"52",
          8607 => x"ff",
          8608 => x"79",
          8609 => x"7b",
          8610 => x"06",
          8611 => x"51",
          8612 => x"3f",
          8613 => x"1c",
          8614 => x"32",
          8615 => x"96",
          8616 => x"06",
          8617 => x"91",
          8618 => x"a1",
          8619 => x"55",
          8620 => x"ff",
          8621 => x"74",
          8622 => x"06",
          8623 => x"51",
          8624 => x"3f",
          8625 => x"52",
          8626 => x"ff",
          8627 => x"f8",
          8628 => x"34",
          8629 => x"1b",
          8630 => x"d9",
          8631 => x"52",
          8632 => x"ff",
          8633 => x"60",
          8634 => x"51",
          8635 => x"3f",
          8636 => x"09",
          8637 => x"cb",
          8638 => x"b2",
          8639 => x"c3",
          8640 => x"a0",
          8641 => x"52",
          8642 => x"ff",
          8643 => x"82",
          8644 => x"51",
          8645 => x"3f",
          8646 => x"1b",
          8647 => x"95",
          8648 => x"b2",
          8649 => x"a0",
          8650 => x"80",
          8651 => x"1c",
          8652 => x"80",
          8653 => x"93",
          8654 => x"a8",
          8655 => x"1b",
          8656 => x"82",
          8657 => x"52",
          8658 => x"ff",
          8659 => x"7c",
          8660 => x"06",
          8661 => x"51",
          8662 => x"3f",
          8663 => x"a4",
          8664 => x"0b",
          8665 => x"93",
          8666 => x"bc",
          8667 => x"51",
          8668 => x"3f",
          8669 => x"52",
          8670 => x"70",
          8671 => x"9f",
          8672 => x"54",
          8673 => x"52",
          8674 => x"9b",
          8675 => x"56",
          8676 => x"08",
          8677 => x"7d",
          8678 => x"81",
          8679 => x"38",
          8680 => x"86",
          8681 => x"52",
          8682 => x"9b",
          8683 => x"80",
          8684 => x"7a",
          8685 => x"ed",
          8686 => x"85",
          8687 => x"7a",
          8688 => x"8f",
          8689 => x"85",
          8690 => x"83",
          8691 => x"ff",
          8692 => x"ff",
          8693 => x"e8",
          8694 => x"9e",
          8695 => x"52",
          8696 => x"51",
          8697 => x"3f",
          8698 => x"52",
          8699 => x"9e",
          8700 => x"54",
          8701 => x"53",
          8702 => x"51",
          8703 => x"3f",
          8704 => x"16",
          8705 => x"7e",
          8706 => x"d8",
          8707 => x"80",
          8708 => x"ff",
          8709 => x"7f",
          8710 => x"7d",
          8711 => x"81",
          8712 => x"f8",
          8713 => x"ff",
          8714 => x"ff",
          8715 => x"51",
          8716 => x"3f",
          8717 => x"88",
          8718 => x"39",
          8719 => x"f8",
          8720 => x"2e",
          8721 => x"55",
          8722 => x"51",
          8723 => x"3f",
          8724 => x"57",
          8725 => x"83",
          8726 => x"76",
          8727 => x"7a",
          8728 => x"ff",
          8729 => x"82",
          8730 => x"82",
          8731 => x"80",
          8732 => x"98",
          8733 => x"51",
          8734 => x"3f",
          8735 => x"78",
          8736 => x"74",
          8737 => x"18",
          8738 => x"2e",
          8739 => x"79",
          8740 => x"2e",
          8741 => x"55",
          8742 => x"62",
          8743 => x"74",
          8744 => x"75",
          8745 => x"7e",
          8746 => x"b8",
          8747 => x"98",
          8748 => x"38",
          8749 => x"78",
          8750 => x"74",
          8751 => x"56",
          8752 => x"93",
          8753 => x"66",
          8754 => x"26",
          8755 => x"56",
          8756 => x"83",
          8757 => x"64",
          8758 => x"77",
          8759 => x"84",
          8760 => x"52",
          8761 => x"9d",
          8762 => x"d4",
          8763 => x"51",
          8764 => x"3f",
          8765 => x"55",
          8766 => x"81",
          8767 => x"34",
          8768 => x"16",
          8769 => x"16",
          8770 => x"16",
          8771 => x"05",
          8772 => x"c1",
          8773 => x"fe",
          8774 => x"fe",
          8775 => x"34",
          8776 => x"08",
          8777 => x"07",
          8778 => x"16",
          8779 => x"98",
          8780 => x"34",
          8781 => x"c6",
          8782 => x"9c",
          8783 => x"52",
          8784 => x"51",
          8785 => x"3f",
          8786 => x"53",
          8787 => x"51",
          8788 => x"3f",
          8789 => x"b6",
          8790 => x"38",
          8791 => x"52",
          8792 => x"99",
          8793 => x"56",
          8794 => x"08",
          8795 => x"39",
          8796 => x"39",
          8797 => x"39",
          8798 => x"08",
          8799 => x"b6",
          8800 => x"3d",
          8801 => x"3d",
          8802 => x"5b",
          8803 => x"60",
          8804 => x"57",
          8805 => x"25",
          8806 => x"3d",
          8807 => x"55",
          8808 => x"15",
          8809 => x"c9",
          8810 => x"81",
          8811 => x"06",
          8812 => x"3d",
          8813 => x"8d",
          8814 => x"74",
          8815 => x"05",
          8816 => x"17",
          8817 => x"2e",
          8818 => x"c9",
          8819 => x"34",
          8820 => x"83",
          8821 => x"74",
          8822 => x"0c",
          8823 => x"04",
          8824 => x"7b",
          8825 => x"b3",
          8826 => x"57",
          8827 => x"09",
          8828 => x"38",
          8829 => x"51",
          8830 => x"17",
          8831 => x"76",
          8832 => x"88",
          8833 => x"17",
          8834 => x"59",
          8835 => x"81",
          8836 => x"76",
          8837 => x"8b",
          8838 => x"54",
          8839 => x"17",
          8840 => x"51",
          8841 => x"79",
          8842 => x"30",
          8843 => x"9f",
          8844 => x"53",
          8845 => x"75",
          8846 => x"81",
          8847 => x"0c",
          8848 => x"04",
          8849 => x"79",
          8850 => x"56",
          8851 => x"24",
          8852 => x"3d",
          8853 => x"74",
          8854 => x"52",
          8855 => x"cb",
          8856 => x"b6",
          8857 => x"38",
          8858 => x"78",
          8859 => x"06",
          8860 => x"16",
          8861 => x"39",
          8862 => x"82",
          8863 => x"89",
          8864 => x"fd",
          8865 => x"54",
          8866 => x"80",
          8867 => x"ff",
          8868 => x"76",
          8869 => x"3d",
          8870 => x"3d",
          8871 => x"e3",
          8872 => x"53",
          8873 => x"53",
          8874 => x"3f",
          8875 => x"51",
          8876 => x"72",
          8877 => x"3f",
          8878 => x"04",
          8879 => x"ff",
          8880 => x"00",
          8881 => x"ff",
          8882 => x"ff",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"69",
          9020 => x"00",
          9021 => x"69",
          9022 => x"6c",
          9023 => x"69",
          9024 => x"00",
          9025 => x"6c",
          9026 => x"00",
          9027 => x"65",
          9028 => x"00",
          9029 => x"63",
          9030 => x"72",
          9031 => x"63",
          9032 => x"00",
          9033 => x"64",
          9034 => x"00",
          9035 => x"64",
          9036 => x"00",
          9037 => x"65",
          9038 => x"65",
          9039 => x"65",
          9040 => x"69",
          9041 => x"69",
          9042 => x"66",
          9043 => x"66",
          9044 => x"61",
          9045 => x"00",
          9046 => x"6d",
          9047 => x"65",
          9048 => x"72",
          9049 => x"65",
          9050 => x"00",
          9051 => x"6e",
          9052 => x"00",
          9053 => x"65",
          9054 => x"00",
          9055 => x"62",
          9056 => x"63",
          9057 => x"62",
          9058 => x"63",
          9059 => x"69",
          9060 => x"00",
          9061 => x"64",
          9062 => x"69",
          9063 => x"45",
          9064 => x"72",
          9065 => x"6e",
          9066 => x"6e",
          9067 => x"65",
          9068 => x"72",
          9069 => x"69",
          9070 => x"6e",
          9071 => x"72",
          9072 => x"79",
          9073 => x"6f",
          9074 => x"6c",
          9075 => x"6f",
          9076 => x"2e",
          9077 => x"6f",
          9078 => x"74",
          9079 => x"6f",
          9080 => x"2e",
          9081 => x"6e",
          9082 => x"69",
          9083 => x"69",
          9084 => x"61",
          9085 => x"00",
          9086 => x"63",
          9087 => x"73",
          9088 => x"6e",
          9089 => x"2e",
          9090 => x"69",
          9091 => x"61",
          9092 => x"61",
          9093 => x"65",
          9094 => x"74",
          9095 => x"00",
          9096 => x"69",
          9097 => x"68",
          9098 => x"6c",
          9099 => x"6e",
          9100 => x"69",
          9101 => x"00",
          9102 => x"44",
          9103 => x"20",
          9104 => x"74",
          9105 => x"72",
          9106 => x"63",
          9107 => x"2e",
          9108 => x"72",
          9109 => x"20",
          9110 => x"62",
          9111 => x"69",
          9112 => x"6e",
          9113 => x"69",
          9114 => x"00",
          9115 => x"69",
          9116 => x"6e",
          9117 => x"65",
          9118 => x"6c",
          9119 => x"00",
          9120 => x"6f",
          9121 => x"6d",
          9122 => x"69",
          9123 => x"20",
          9124 => x"65",
          9125 => x"74",
          9126 => x"66",
          9127 => x"64",
          9128 => x"20",
          9129 => x"6b",
          9130 => x"6f",
          9131 => x"74",
          9132 => x"6f",
          9133 => x"64",
          9134 => x"69",
          9135 => x"75",
          9136 => x"6f",
          9137 => x"61",
          9138 => x"6e",
          9139 => x"6e",
          9140 => x"6c",
          9141 => x"00",
          9142 => x"69",
          9143 => x"69",
          9144 => x"6f",
          9145 => x"64",
          9146 => x"6e",
          9147 => x"66",
          9148 => x"65",
          9149 => x"6d",
          9150 => x"72",
          9151 => x"00",
          9152 => x"6f",
          9153 => x"61",
          9154 => x"6f",
          9155 => x"20",
          9156 => x"65",
          9157 => x"00",
          9158 => x"61",
          9159 => x"65",
          9160 => x"73",
          9161 => x"63",
          9162 => x"65",
          9163 => x"00",
          9164 => x"75",
          9165 => x"73",
          9166 => x"00",
          9167 => x"6e",
          9168 => x"77",
          9169 => x"72",
          9170 => x"2e",
          9171 => x"25",
          9172 => x"62",
          9173 => x"73",
          9174 => x"20",
          9175 => x"25",
          9176 => x"62",
          9177 => x"73",
          9178 => x"63",
          9179 => x"00",
          9180 => x"65",
          9181 => x"00",
          9182 => x"3d",
          9183 => x"6c",
          9184 => x"31",
          9185 => x"38",
          9186 => x"20",
          9187 => x"30",
          9188 => x"2c",
          9189 => x"4f",
          9190 => x"30",
          9191 => x"20",
          9192 => x"6c",
          9193 => x"30",
          9194 => x"0a",
          9195 => x"30",
          9196 => x"00",
          9197 => x"20",
          9198 => x"30",
          9199 => x"00",
          9200 => x"20",
          9201 => x"20",
          9202 => x"00",
          9203 => x"30",
          9204 => x"00",
          9205 => x"20",
          9206 => x"7c",
          9207 => x"00",
          9208 => x"4f",
          9209 => x"2a",
          9210 => x"73",
          9211 => x"00",
          9212 => x"32",
          9213 => x"2f",
          9214 => x"30",
          9215 => x"31",
          9216 => x"00",
          9217 => x"5a",
          9218 => x"20",
          9219 => x"20",
          9220 => x"78",
          9221 => x"73",
          9222 => x"20",
          9223 => x"0a",
          9224 => x"50",
          9225 => x"6e",
          9226 => x"72",
          9227 => x"20",
          9228 => x"64",
          9229 => x"00",
          9230 => x"69",
          9231 => x"20",
          9232 => x"65",
          9233 => x"70",
          9234 => x"53",
          9235 => x"6e",
          9236 => x"72",
          9237 => x"00",
          9238 => x"4f",
          9239 => x"20",
          9240 => x"69",
          9241 => x"72",
          9242 => x"74",
          9243 => x"4f",
          9244 => x"20",
          9245 => x"69",
          9246 => x"72",
          9247 => x"74",
          9248 => x"41",
          9249 => x"20",
          9250 => x"69",
          9251 => x"72",
          9252 => x"74",
          9253 => x"41",
          9254 => x"20",
          9255 => x"69",
          9256 => x"72",
          9257 => x"74",
          9258 => x"41",
          9259 => x"20",
          9260 => x"69",
          9261 => x"72",
          9262 => x"74",
          9263 => x"41",
          9264 => x"20",
          9265 => x"69",
          9266 => x"72",
          9267 => x"74",
          9268 => x"65",
          9269 => x"6e",
          9270 => x"70",
          9271 => x"6d",
          9272 => x"2e",
          9273 => x"6e",
          9274 => x"69",
          9275 => x"74",
          9276 => x"72",
          9277 => x"00",
          9278 => x"75",
          9279 => x"78",
          9280 => x"62",
          9281 => x"00",
          9282 => x"4f",
          9283 => x"73",
          9284 => x"3a",
          9285 => x"61",
          9286 => x"64",
          9287 => x"20",
          9288 => x"74",
          9289 => x"69",
          9290 => x"73",
          9291 => x"61",
          9292 => x"30",
          9293 => x"6c",
          9294 => x"65",
          9295 => x"69",
          9296 => x"61",
          9297 => x"6c",
          9298 => x"00",
          9299 => x"20",
          9300 => x"6c",
          9301 => x"69",
          9302 => x"2e",
          9303 => x"00",
          9304 => x"6f",
          9305 => x"6e",
          9306 => x"2e",
          9307 => x"6f",
          9308 => x"72",
          9309 => x"2e",
          9310 => x"00",
          9311 => x"30",
          9312 => x"28",
          9313 => x"78",
          9314 => x"25",
          9315 => x"78",
          9316 => x"38",
          9317 => x"00",
          9318 => x"75",
          9319 => x"4d",
          9320 => x"72",
          9321 => x"43",
          9322 => x"6c",
          9323 => x"2e",
          9324 => x"30",
          9325 => x"20",
          9326 => x"58",
          9327 => x"3f",
          9328 => x"30",
          9329 => x"20",
          9330 => x"58",
          9331 => x"30",
          9332 => x"20",
          9333 => x"6c",
          9334 => x"00",
          9335 => x"78",
          9336 => x"74",
          9337 => x"20",
          9338 => x"65",
          9339 => x"25",
          9340 => x"78",
          9341 => x"2e",
          9342 => x"61",
          9343 => x"6e",
          9344 => x"6f",
          9345 => x"40",
          9346 => x"38",
          9347 => x"2e",
          9348 => x"00",
          9349 => x"61",
          9350 => x"72",
          9351 => x"72",
          9352 => x"20",
          9353 => x"65",
          9354 => x"64",
          9355 => x"00",
          9356 => x"65",
          9357 => x"72",
          9358 => x"67",
          9359 => x"70",
          9360 => x"61",
          9361 => x"6e",
          9362 => x"00",
          9363 => x"6f",
          9364 => x"72",
          9365 => x"6f",
          9366 => x"67",
          9367 => x"00",
          9368 => x"50",
          9369 => x"69",
          9370 => x"64",
          9371 => x"73",
          9372 => x"2e",
          9373 => x"00",
          9374 => x"64",
          9375 => x"73",
          9376 => x"00",
          9377 => x"64",
          9378 => x"73",
          9379 => x"61",
          9380 => x"6f",
          9381 => x"6e",
          9382 => x"00",
          9383 => x"75",
          9384 => x"6e",
          9385 => x"2e",
          9386 => x"6e",
          9387 => x"69",
          9388 => x"69",
          9389 => x"72",
          9390 => x"74",
          9391 => x"2e",
          9392 => x"64",
          9393 => x"2f",
          9394 => x"25",
          9395 => x"64",
          9396 => x"2e",
          9397 => x"64",
          9398 => x"6f",
          9399 => x"6f",
          9400 => x"67",
          9401 => x"74",
          9402 => x"00",
          9403 => x"28",
          9404 => x"6d",
          9405 => x"43",
          9406 => x"6e",
          9407 => x"29",
          9408 => x"0a",
          9409 => x"69",
          9410 => x"20",
          9411 => x"6c",
          9412 => x"6e",
          9413 => x"3a",
          9414 => x"20",
          9415 => x"42",
          9416 => x"52",
          9417 => x"20",
          9418 => x"38",
          9419 => x"30",
          9420 => x"2e",
          9421 => x"20",
          9422 => x"44",
          9423 => x"20",
          9424 => x"20",
          9425 => x"38",
          9426 => x"30",
          9427 => x"2e",
          9428 => x"20",
          9429 => x"4e",
          9430 => x"42",
          9431 => x"20",
          9432 => x"38",
          9433 => x"30",
          9434 => x"2e",
          9435 => x"20",
          9436 => x"52",
          9437 => x"20",
          9438 => x"20",
          9439 => x"38",
          9440 => x"30",
          9441 => x"2e",
          9442 => x"20",
          9443 => x"41",
          9444 => x"20",
          9445 => x"20",
          9446 => x"38",
          9447 => x"30",
          9448 => x"2e",
          9449 => x"20",
          9450 => x"44",
          9451 => x"52",
          9452 => x"20",
          9453 => x"76",
          9454 => x"73",
          9455 => x"30",
          9456 => x"2e",
          9457 => x"20",
          9458 => x"49",
          9459 => x"31",
          9460 => x"20",
          9461 => x"6d",
          9462 => x"20",
          9463 => x"30",
          9464 => x"2e",
          9465 => x"20",
          9466 => x"4e",
          9467 => x"43",
          9468 => x"20",
          9469 => x"61",
          9470 => x"6c",
          9471 => x"30",
          9472 => x"2e",
          9473 => x"20",
          9474 => x"49",
          9475 => x"4f",
          9476 => x"42",
          9477 => x"00",
          9478 => x"20",
          9479 => x"42",
          9480 => x"43",
          9481 => x"20",
          9482 => x"4f",
          9483 => x"00",
          9484 => x"20",
          9485 => x"53",
          9486 => x"20",
          9487 => x"50",
          9488 => x"64",
          9489 => x"73",
          9490 => x"3a",
          9491 => x"20",
          9492 => x"50",
          9493 => x"65",
          9494 => x"20",
          9495 => x"74",
          9496 => x"41",
          9497 => x"65",
          9498 => x"3d",
          9499 => x"38",
          9500 => x"00",
          9501 => x"20",
          9502 => x"50",
          9503 => x"65",
          9504 => x"79",
          9505 => x"61",
          9506 => x"41",
          9507 => x"65",
          9508 => x"3d",
          9509 => x"38",
          9510 => x"00",
          9511 => x"20",
          9512 => x"74",
          9513 => x"20",
          9514 => x"72",
          9515 => x"64",
          9516 => x"73",
          9517 => x"20",
          9518 => x"3d",
          9519 => x"38",
          9520 => x"00",
          9521 => x"69",
          9522 => x"00",
          9523 => x"20",
          9524 => x"50",
          9525 => x"64",
          9526 => x"20",
          9527 => x"20",
          9528 => x"20",
          9529 => x"20",
          9530 => x"3d",
          9531 => x"34",
          9532 => x"00",
          9533 => x"20",
          9534 => x"79",
          9535 => x"6d",
          9536 => x"6f",
          9537 => x"46",
          9538 => x"20",
          9539 => x"20",
          9540 => x"3d",
          9541 => x"2e",
          9542 => x"64",
          9543 => x"0a",
          9544 => x"20",
          9545 => x"44",
          9546 => x"20",
          9547 => x"63",
          9548 => x"72",
          9549 => x"20",
          9550 => x"20",
          9551 => x"3d",
          9552 => x"2e",
          9553 => x"64",
          9554 => x"0a",
          9555 => x"20",
          9556 => x"69",
          9557 => x"6f",
          9558 => x"53",
          9559 => x"4d",
          9560 => x"6f",
          9561 => x"46",
          9562 => x"3d",
          9563 => x"2e",
          9564 => x"64",
          9565 => x"0a",
          9566 => x"6d",
          9567 => x"00",
          9568 => x"65",
          9569 => x"6d",
          9570 => x"6c",
          9571 => x"00",
          9572 => x"56",
          9573 => x"56",
          9574 => x"00",
          9575 => x"6e",
          9576 => x"77",
          9577 => x"00",
          9578 => x"00",
          9579 => x"00",
          9580 => x"00",
          9581 => x"00",
          9582 => x"00",
          9583 => x"00",
          9584 => x"00",
          9585 => x"00",
          9586 => x"00",
          9587 => x"00",
          9588 => x"00",
          9589 => x"00",
          9590 => x"00",
          9591 => x"00",
          9592 => x"00",
          9593 => x"00",
          9594 => x"00",
          9595 => x"00",
          9596 => x"00",
          9597 => x"00",
          9598 => x"00",
          9599 => x"00",
          9600 => x"00",
          9601 => x"00",
          9602 => x"00",
          9603 => x"00",
          9604 => x"00",
          9605 => x"00",
          9606 => x"00",
          9607 => x"00",
          9608 => x"00",
          9609 => x"00",
          9610 => x"00",
          9611 => x"00",
          9612 => x"00",
          9613 => x"00",
          9614 => x"00",
          9615 => x"00",
          9616 => x"00",
          9617 => x"00",
          9618 => x"00",
          9619 => x"00",
          9620 => x"00",
          9621 => x"00",
          9622 => x"00",
          9623 => x"00",
          9624 => x"00",
          9625 => x"00",
          9626 => x"00",
          9627 => x"00",
          9628 => x"00",
          9629 => x"00",
          9630 => x"00",
          9631 => x"00",
          9632 => x"00",
          9633 => x"00",
          9634 => x"00",
          9635 => x"00",
          9636 => x"00",
          9637 => x"00",
          9638 => x"00",
          9639 => x"00",
          9640 => x"00",
          9641 => x"00",
          9642 => x"00",
          9643 => x"5b",
          9644 => x"5b",
          9645 => x"5b",
          9646 => x"5b",
          9647 => x"5b",
          9648 => x"5b",
          9649 => x"5b",
          9650 => x"30",
          9651 => x"5b",
          9652 => x"5b",
          9653 => x"5b",
          9654 => x"00",
          9655 => x"00",
          9656 => x"00",
          9657 => x"00",
          9658 => x"00",
          9659 => x"00",
          9660 => x"00",
          9661 => x"00",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"69",
          9666 => x"72",
          9667 => x"69",
          9668 => x"00",
          9669 => x"00",
          9670 => x"30",
          9671 => x"20",
          9672 => x"0a",
          9673 => x"61",
          9674 => x"64",
          9675 => x"20",
          9676 => x"65",
          9677 => x"68",
          9678 => x"69",
          9679 => x"72",
          9680 => x"69",
          9681 => x"74",
          9682 => x"4f",
          9683 => x"00",
          9684 => x"61",
          9685 => x"74",
          9686 => x"65",
          9687 => x"72",
          9688 => x"65",
          9689 => x"73",
          9690 => x"79",
          9691 => x"6c",
          9692 => x"64",
          9693 => x"62",
          9694 => x"67",
          9695 => x"44",
          9696 => x"2a",
          9697 => x"3b",
          9698 => x"3f",
          9699 => x"7f",
          9700 => x"41",
          9701 => x"41",
          9702 => x"00",
          9703 => x"fe",
          9704 => x"44",
          9705 => x"2e",
          9706 => x"4f",
          9707 => x"4d",
          9708 => x"20",
          9709 => x"54",
          9710 => x"20",
          9711 => x"4f",
          9712 => x"4d",
          9713 => x"20",
          9714 => x"54",
          9715 => x"20",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"9a",
          9721 => x"41",
          9722 => x"45",
          9723 => x"49",
          9724 => x"92",
          9725 => x"4f",
          9726 => x"99",
          9727 => x"9d",
          9728 => x"49",
          9729 => x"a5",
          9730 => x"a9",
          9731 => x"ad",
          9732 => x"b1",
          9733 => x"b5",
          9734 => x"b9",
          9735 => x"bd",
          9736 => x"c1",
          9737 => x"c5",
          9738 => x"c9",
          9739 => x"cd",
          9740 => x"d1",
          9741 => x"d5",
          9742 => x"d9",
          9743 => x"dd",
          9744 => x"e1",
          9745 => x"e5",
          9746 => x"e9",
          9747 => x"ed",
          9748 => x"f1",
          9749 => x"f5",
          9750 => x"f9",
          9751 => x"fd",
          9752 => x"2e",
          9753 => x"5b",
          9754 => x"22",
          9755 => x"3e",
          9756 => x"00",
          9757 => x"01",
          9758 => x"10",
          9759 => x"00",
          9760 => x"00",
          9761 => x"01",
          9762 => x"04",
          9763 => x"10",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"02",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"04",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"14",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"2b",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"30",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"3c",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"3d",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"3f",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"40",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"41",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"42",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"43",
          9812 => x"00",
          9813 => x"00",
          9814 => x"00",
          9815 => x"50",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"51",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"54",
          9824 => x"00",
          9825 => x"00",
          9826 => x"00",
          9827 => x"55",
          9828 => x"00",
          9829 => x"00",
          9830 => x"00",
          9831 => x"79",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"78",
          9836 => x"00",
          9837 => x"00",
          9838 => x"00",
          9839 => x"82",
          9840 => x"00",
          9841 => x"00",
          9842 => x"00",
          9843 => x"83",
          9844 => x"00",
          9845 => x"00",
          9846 => x"00",
          9847 => x"85",
          9848 => x"00",
          9849 => x"00",
          9850 => x"00",
          9851 => x"87",
          9852 => x"00",
          9853 => x"00",
          9854 => x"00",
          9855 => x"8c",
          9856 => x"00",
          9857 => x"00",
          9858 => x"00",
          9859 => x"8d",
          9860 => x"00",
          9861 => x"00",
          9862 => x"00",
          9863 => x"8e",
          9864 => x"00",
          9865 => x"00",
          9866 => x"00",
          9867 => x"8f",
          9868 => x"00",
          9869 => x"00",
          9870 => x"00",
          9871 => x"00",
          9872 => x"00",
          9873 => x"00",
          9874 => x"00",
          9875 => x"01",
          9876 => x"00",
          9877 => x"01",
          9878 => x"81",
          9879 => x"00",
          9880 => x"7f",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"f5",
          9886 => x"f5",
          9887 => x"f5",
          9888 => x"00",
          9889 => x"01",
          9890 => x"01",
          9891 => x"01",
          9892 => x"00",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"00",
          9898 => x"00",
          9899 => x"00",
          9900 => x"00",
          9901 => x"00",
          9902 => x"00",
          9903 => x"00",
          9904 => x"00",
          9905 => x"00",
          9906 => x"00",
          9907 => x"00",
          9908 => x"00",
          9909 => x"00",
          9910 => x"00",
          9911 => x"00",
          9912 => x"00",
          9913 => x"00",
          9914 => x"00",
          9915 => x"00",
          9916 => x"00",
          9917 => x"00",
          9918 => x"00",
          9919 => x"00",
          9920 => x"00",
          9921 => x"00",
          9922 => x"00",
          9923 => x"00",
          9924 => x"00",
          9925 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"9d",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"bc",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"f4",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"e0",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b3",
           272 => x"0b",
           273 => x"0b",
           274 => x"d1",
           275 => x"0b",
           276 => x"0b",
           277 => x"f0",
           278 => x"0b",
           279 => x"0b",
           280 => x"8f",
           281 => x"0b",
           282 => x"0b",
           283 => x"ad",
           284 => x"0b",
           285 => x"0b",
           286 => x"cd",
           287 => x"0b",
           288 => x"0b",
           289 => x"ed",
           290 => x"0b",
           291 => x"0b",
           292 => x"8d",
           293 => x"0b",
           294 => x"0b",
           295 => x"ad",
           296 => x"0b",
           297 => x"0b",
           298 => x"cd",
           299 => x"0b",
           300 => x"0b",
           301 => x"ed",
           302 => x"0b",
           303 => x"0b",
           304 => x"8d",
           305 => x"0b",
           306 => x"0b",
           307 => x"ad",
           308 => x"0b",
           309 => x"0b",
           310 => x"cd",
           311 => x"0b",
           312 => x"0b",
           313 => x"ed",
           314 => x"0b",
           315 => x"0b",
           316 => x"8d",
           317 => x"0b",
           318 => x"0b",
           319 => x"ad",
           320 => x"0b",
           321 => x"0b",
           322 => x"cd",
           323 => x"0b",
           324 => x"0b",
           325 => x"ed",
           326 => x"0b",
           327 => x"0b",
           328 => x"8d",
           329 => x"0b",
           330 => x"0b",
           331 => x"ad",
           332 => x"0b",
           333 => x"0b",
           334 => x"cd",
           335 => x"0b",
           336 => x"0b",
           337 => x"ed",
           338 => x"0b",
           339 => x"0b",
           340 => x"8d",
           341 => x"0b",
           342 => x"0b",
           343 => x"ad",
           344 => x"0b",
           345 => x"0b",
           346 => x"cd",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"82",
           393 => x"82",
           394 => x"af",
           395 => x"b6",
           396 => x"d0",
           397 => x"b6",
           398 => x"ad",
           399 => x"a4",
           400 => x"90",
           401 => x"a4",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"82",
           407 => x"82",
           408 => x"82",
           409 => x"80",
           410 => x"82",
           411 => x"82",
           412 => x"82",
           413 => x"80",
           414 => x"82",
           415 => x"82",
           416 => x"82",
           417 => x"93",
           418 => x"b6",
           419 => x"d0",
           420 => x"b6",
           421 => x"c0",
           422 => x"a4",
           423 => x"90",
           424 => x"a4",
           425 => x"2d",
           426 => x"08",
           427 => x"04",
           428 => x"0c",
           429 => x"2d",
           430 => x"08",
           431 => x"04",
           432 => x"0c",
           433 => x"2d",
           434 => x"08",
           435 => x"04",
           436 => x"0c",
           437 => x"2d",
           438 => x"08",
           439 => x"04",
           440 => x"0c",
           441 => x"2d",
           442 => x"08",
           443 => x"04",
           444 => x"0c",
           445 => x"2d",
           446 => x"08",
           447 => x"04",
           448 => x"0c",
           449 => x"2d",
           450 => x"08",
           451 => x"04",
           452 => x"0c",
           453 => x"2d",
           454 => x"08",
           455 => x"04",
           456 => x"0c",
           457 => x"2d",
           458 => x"08",
           459 => x"04",
           460 => x"0c",
           461 => x"2d",
           462 => x"08",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"04",
           480 => x"0c",
           481 => x"2d",
           482 => x"08",
           483 => x"04",
           484 => x"0c",
           485 => x"2d",
           486 => x"08",
           487 => x"04",
           488 => x"0c",
           489 => x"2d",
           490 => x"08",
           491 => x"04",
           492 => x"0c",
           493 => x"2d",
           494 => x"08",
           495 => x"04",
           496 => x"0c",
           497 => x"2d",
           498 => x"08",
           499 => x"04",
           500 => x"0c",
           501 => x"2d",
           502 => x"08",
           503 => x"04",
           504 => x"0c",
           505 => x"2d",
           506 => x"08",
           507 => x"04",
           508 => x"0c",
           509 => x"2d",
           510 => x"08",
           511 => x"04",
           512 => x"0c",
           513 => x"2d",
           514 => x"08",
           515 => x"04",
           516 => x"0c",
           517 => x"2d",
           518 => x"08",
           519 => x"04",
           520 => x"0c",
           521 => x"2d",
           522 => x"08",
           523 => x"04",
           524 => x"0c",
           525 => x"2d",
           526 => x"08",
           527 => x"04",
           528 => x"0c",
           529 => x"2d",
           530 => x"08",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"04",
           548 => x"0c",
           549 => x"2d",
           550 => x"08",
           551 => x"04",
           552 => x"0c",
           553 => x"2d",
           554 => x"08",
           555 => x"04",
           556 => x"0c",
           557 => x"2d",
           558 => x"08",
           559 => x"04",
           560 => x"0c",
           561 => x"2d",
           562 => x"08",
           563 => x"04",
           564 => x"0c",
           565 => x"2d",
           566 => x"08",
           567 => x"04",
           568 => x"0c",
           569 => x"2d",
           570 => x"08",
           571 => x"04",
           572 => x"0c",
           573 => x"2d",
           574 => x"08",
           575 => x"04",
           576 => x"0c",
           577 => x"2d",
           578 => x"08",
           579 => x"04",
           580 => x"0c",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"0c",
           589 => x"2d",
           590 => x"08",
           591 => x"04",
           592 => x"0c",
           593 => x"2d",
           594 => x"08",
           595 => x"04",
           596 => x"0c",
           597 => x"2d",
           598 => x"08",
           599 => x"04",
           600 => x"00",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"53",
           609 => x"00",
           610 => x"06",
           611 => x"09",
           612 => x"05",
           613 => x"2b",
           614 => x"06",
           615 => x"04",
           616 => x"72",
           617 => x"05",
           618 => x"05",
           619 => x"72",
           620 => x"53",
           621 => x"51",
           622 => x"04",
           623 => x"70",
           624 => x"27",
           625 => x"71",
           626 => x"53",
           627 => x"0b",
           628 => x"8c",
           629 => x"ef",
           630 => x"82",
           631 => x"02",
           632 => x"0c",
           633 => x"82",
           634 => x"8c",
           635 => x"b6",
           636 => x"05",
           637 => x"a4",
           638 => x"08",
           639 => x"a4",
           640 => x"08",
           641 => x"ec",
           642 => x"84",
           643 => x"b6",
           644 => x"82",
           645 => x"f8",
           646 => x"b6",
           647 => x"05",
           648 => x"b6",
           649 => x"54",
           650 => x"82",
           651 => x"04",
           652 => x"08",
           653 => x"a4",
           654 => x"0d",
           655 => x"08",
           656 => x"85",
           657 => x"81",
           658 => x"06",
           659 => x"52",
           660 => x"80",
           661 => x"a4",
           662 => x"08",
           663 => x"8d",
           664 => x"82",
           665 => x"f4",
           666 => x"c4",
           667 => x"a4",
           668 => x"08",
           669 => x"b6",
           670 => x"05",
           671 => x"82",
           672 => x"f8",
           673 => x"b6",
           674 => x"05",
           675 => x"a4",
           676 => x"0c",
           677 => x"08",
           678 => x"8a",
           679 => x"38",
           680 => x"b6",
           681 => x"05",
           682 => x"e9",
           683 => x"a4",
           684 => x"08",
           685 => x"3f",
           686 => x"08",
           687 => x"a4",
           688 => x"0c",
           689 => x"a4",
           690 => x"08",
           691 => x"81",
           692 => x"80",
           693 => x"a4",
           694 => x"0c",
           695 => x"82",
           696 => x"fc",
           697 => x"b6",
           698 => x"05",
           699 => x"71",
           700 => x"b6",
           701 => x"05",
           702 => x"82",
           703 => x"8c",
           704 => x"b6",
           705 => x"05",
           706 => x"82",
           707 => x"fc",
           708 => x"80",
           709 => x"a4",
           710 => x"08",
           711 => x"34",
           712 => x"08",
           713 => x"70",
           714 => x"08",
           715 => x"52",
           716 => x"08",
           717 => x"82",
           718 => x"87",
           719 => x"b6",
           720 => x"82",
           721 => x"02",
           722 => x"0c",
           723 => x"86",
           724 => x"a4",
           725 => x"34",
           726 => x"08",
           727 => x"82",
           728 => x"e0",
           729 => x"0a",
           730 => x"a4",
           731 => x"0c",
           732 => x"08",
           733 => x"82",
           734 => x"fc",
           735 => x"b6",
           736 => x"05",
           737 => x"b6",
           738 => x"05",
           739 => x"b6",
           740 => x"05",
           741 => x"54",
           742 => x"82",
           743 => x"70",
           744 => x"08",
           745 => x"82",
           746 => x"ec",
           747 => x"b6",
           748 => x"05",
           749 => x"54",
           750 => x"82",
           751 => x"dc",
           752 => x"82",
           753 => x"54",
           754 => x"82",
           755 => x"04",
           756 => x"08",
           757 => x"a4",
           758 => x"0d",
           759 => x"08",
           760 => x"82",
           761 => x"fc",
           762 => x"b6",
           763 => x"05",
           764 => x"b6",
           765 => x"05",
           766 => x"b6",
           767 => x"05",
           768 => x"a3",
           769 => x"98",
           770 => x"b6",
           771 => x"05",
           772 => x"a4",
           773 => x"08",
           774 => x"98",
           775 => x"87",
           776 => x"b6",
           777 => x"82",
           778 => x"02",
           779 => x"0c",
           780 => x"80",
           781 => x"a4",
           782 => x"23",
           783 => x"08",
           784 => x"53",
           785 => x"14",
           786 => x"a4",
           787 => x"08",
           788 => x"70",
           789 => x"81",
           790 => x"06",
           791 => x"51",
           792 => x"2e",
           793 => x"0b",
           794 => x"08",
           795 => x"96",
           796 => x"b6",
           797 => x"05",
           798 => x"33",
           799 => x"b6",
           800 => x"05",
           801 => x"ff",
           802 => x"80",
           803 => x"38",
           804 => x"08",
           805 => x"81",
           806 => x"a4",
           807 => x"0c",
           808 => x"08",
           809 => x"70",
           810 => x"53",
           811 => x"95",
           812 => x"b6",
           813 => x"05",
           814 => x"73",
           815 => x"38",
           816 => x"08",
           817 => x"53",
           818 => x"81",
           819 => x"b6",
           820 => x"05",
           821 => x"b0",
           822 => x"06",
           823 => x"82",
           824 => x"e8",
           825 => x"98",
           826 => x"2c",
           827 => x"72",
           828 => x"b6",
           829 => x"05",
           830 => x"2a",
           831 => x"70",
           832 => x"51",
           833 => x"80",
           834 => x"82",
           835 => x"e4",
           836 => x"82",
           837 => x"53",
           838 => x"a4",
           839 => x"23",
           840 => x"82",
           841 => x"e8",
           842 => x"98",
           843 => x"2c",
           844 => x"2b",
           845 => x"11",
           846 => x"53",
           847 => x"72",
           848 => x"08",
           849 => x"82",
           850 => x"e8",
           851 => x"82",
           852 => x"f8",
           853 => x"15",
           854 => x"51",
           855 => x"b6",
           856 => x"05",
           857 => x"a4",
           858 => x"33",
           859 => x"70",
           860 => x"51",
           861 => x"25",
           862 => x"ff",
           863 => x"a4",
           864 => x"34",
           865 => x"08",
           866 => x"70",
           867 => x"81",
           868 => x"53",
           869 => x"38",
           870 => x"08",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"53",
           876 => x"a4",
           877 => x"23",
           878 => x"82",
           879 => x"e4",
           880 => x"83",
           881 => x"06",
           882 => x"72",
           883 => x"38",
           884 => x"08",
           885 => x"70",
           886 => x"98",
           887 => x"53",
           888 => x"81",
           889 => x"a4",
           890 => x"34",
           891 => x"08",
           892 => x"e0",
           893 => x"a4",
           894 => x"0c",
           895 => x"a4",
           896 => x"08",
           897 => x"92",
           898 => x"b6",
           899 => x"05",
           900 => x"2b",
           901 => x"11",
           902 => x"51",
           903 => x"04",
           904 => x"08",
           905 => x"70",
           906 => x"53",
           907 => x"a4",
           908 => x"23",
           909 => x"08",
           910 => x"70",
           911 => x"53",
           912 => x"a4",
           913 => x"23",
           914 => x"82",
           915 => x"e4",
           916 => x"81",
           917 => x"53",
           918 => x"a4",
           919 => x"23",
           920 => x"82",
           921 => x"e4",
           922 => x"80",
           923 => x"53",
           924 => x"a4",
           925 => x"23",
           926 => x"82",
           927 => x"e4",
           928 => x"88",
           929 => x"72",
           930 => x"08",
           931 => x"80",
           932 => x"a4",
           933 => x"34",
           934 => x"82",
           935 => x"e4",
           936 => x"84",
           937 => x"72",
           938 => x"08",
           939 => x"fb",
           940 => x"0b",
           941 => x"08",
           942 => x"82",
           943 => x"ec",
           944 => x"11",
           945 => x"82",
           946 => x"ec",
           947 => x"e3",
           948 => x"a4",
           949 => x"34",
           950 => x"82",
           951 => x"90",
           952 => x"b6",
           953 => x"05",
           954 => x"82",
           955 => x"90",
           956 => x"08",
           957 => x"82",
           958 => x"fc",
           959 => x"b6",
           960 => x"05",
           961 => x"51",
           962 => x"b6",
           963 => x"05",
           964 => x"39",
           965 => x"08",
           966 => x"82",
           967 => x"90",
           968 => x"05",
           969 => x"08",
           970 => x"70",
           971 => x"a4",
           972 => x"0c",
           973 => x"08",
           974 => x"70",
           975 => x"81",
           976 => x"51",
           977 => x"2e",
           978 => x"b6",
           979 => x"05",
           980 => x"2b",
           981 => x"2c",
           982 => x"a4",
           983 => x"08",
           984 => x"d8",
           985 => x"98",
           986 => x"82",
           987 => x"f4",
           988 => x"39",
           989 => x"08",
           990 => x"51",
           991 => x"82",
           992 => x"53",
           993 => x"a4",
           994 => x"23",
           995 => x"08",
           996 => x"53",
           997 => x"08",
           998 => x"73",
           999 => x"54",
          1000 => x"a4",
          1001 => x"23",
          1002 => x"82",
          1003 => x"90",
          1004 => x"b6",
          1005 => x"05",
          1006 => x"82",
          1007 => x"90",
          1008 => x"08",
          1009 => x"08",
          1010 => x"82",
          1011 => x"e4",
          1012 => x"83",
          1013 => x"06",
          1014 => x"53",
          1015 => x"ab",
          1016 => x"a4",
          1017 => x"33",
          1018 => x"53",
          1019 => x"53",
          1020 => x"08",
          1021 => x"52",
          1022 => x"3f",
          1023 => x"08",
          1024 => x"b6",
          1025 => x"05",
          1026 => x"82",
          1027 => x"fc",
          1028 => x"9b",
          1029 => x"b6",
          1030 => x"72",
          1031 => x"08",
          1032 => x"82",
          1033 => x"ec",
          1034 => x"82",
          1035 => x"f4",
          1036 => x"71",
          1037 => x"72",
          1038 => x"08",
          1039 => x"8a",
          1040 => x"b6",
          1041 => x"05",
          1042 => x"2a",
          1043 => x"51",
          1044 => x"80",
          1045 => x"82",
          1046 => x"90",
          1047 => x"b6",
          1048 => x"05",
          1049 => x"82",
          1050 => x"90",
          1051 => x"08",
          1052 => x"08",
          1053 => x"53",
          1054 => x"b6",
          1055 => x"05",
          1056 => x"a4",
          1057 => x"08",
          1058 => x"b6",
          1059 => x"05",
          1060 => x"82",
          1061 => x"dc",
          1062 => x"82",
          1063 => x"dc",
          1064 => x"b6",
          1065 => x"05",
          1066 => x"a4",
          1067 => x"08",
          1068 => x"38",
          1069 => x"08",
          1070 => x"70",
          1071 => x"53",
          1072 => x"a4",
          1073 => x"23",
          1074 => x"08",
          1075 => x"30",
          1076 => x"08",
          1077 => x"82",
          1078 => x"e4",
          1079 => x"ff",
          1080 => x"53",
          1081 => x"a4",
          1082 => x"23",
          1083 => x"88",
          1084 => x"a4",
          1085 => x"23",
          1086 => x"b6",
          1087 => x"05",
          1088 => x"c0",
          1089 => x"72",
          1090 => x"08",
          1091 => x"80",
          1092 => x"b6",
          1093 => x"05",
          1094 => x"82",
          1095 => x"f4",
          1096 => x"b6",
          1097 => x"05",
          1098 => x"2a",
          1099 => x"51",
          1100 => x"80",
          1101 => x"82",
          1102 => x"90",
          1103 => x"b6",
          1104 => x"05",
          1105 => x"82",
          1106 => x"90",
          1107 => x"08",
          1108 => x"08",
          1109 => x"53",
          1110 => x"b6",
          1111 => x"05",
          1112 => x"a4",
          1113 => x"08",
          1114 => x"b6",
          1115 => x"05",
          1116 => x"82",
          1117 => x"d8",
          1118 => x"82",
          1119 => x"d8",
          1120 => x"b6",
          1121 => x"05",
          1122 => x"a4",
          1123 => x"22",
          1124 => x"51",
          1125 => x"b6",
          1126 => x"05",
          1127 => x"a8",
          1128 => x"a4",
          1129 => x"0c",
          1130 => x"08",
          1131 => x"82",
          1132 => x"f4",
          1133 => x"b6",
          1134 => x"05",
          1135 => x"70",
          1136 => x"55",
          1137 => x"82",
          1138 => x"53",
          1139 => x"82",
          1140 => x"f0",
          1141 => x"b6",
          1142 => x"05",
          1143 => x"a4",
          1144 => x"08",
          1145 => x"53",
          1146 => x"a4",
          1147 => x"a4",
          1148 => x"08",
          1149 => x"54",
          1150 => x"08",
          1151 => x"70",
          1152 => x"51",
          1153 => x"82",
          1154 => x"d0",
          1155 => x"39",
          1156 => x"08",
          1157 => x"53",
          1158 => x"11",
          1159 => x"82",
          1160 => x"d0",
          1161 => x"b6",
          1162 => x"05",
          1163 => x"b6",
          1164 => x"05",
          1165 => x"82",
          1166 => x"f0",
          1167 => x"05",
          1168 => x"08",
          1169 => x"82",
          1170 => x"f4",
          1171 => x"53",
          1172 => x"08",
          1173 => x"52",
          1174 => x"3f",
          1175 => x"08",
          1176 => x"a4",
          1177 => x"0c",
          1178 => x"a4",
          1179 => x"08",
          1180 => x"38",
          1181 => x"82",
          1182 => x"f0",
          1183 => x"b6",
          1184 => x"72",
          1185 => x"75",
          1186 => x"72",
          1187 => x"08",
          1188 => x"82",
          1189 => x"e4",
          1190 => x"b2",
          1191 => x"72",
          1192 => x"38",
          1193 => x"08",
          1194 => x"ff",
          1195 => x"72",
          1196 => x"08",
          1197 => x"82",
          1198 => x"e4",
          1199 => x"86",
          1200 => x"06",
          1201 => x"72",
          1202 => x"e7",
          1203 => x"a4",
          1204 => x"22",
          1205 => x"82",
          1206 => x"cc",
          1207 => x"b6",
          1208 => x"05",
          1209 => x"82",
          1210 => x"cc",
          1211 => x"b6",
          1212 => x"05",
          1213 => x"72",
          1214 => x"81",
          1215 => x"82",
          1216 => x"cc",
          1217 => x"05",
          1218 => x"b6",
          1219 => x"05",
          1220 => x"82",
          1221 => x"cc",
          1222 => x"05",
          1223 => x"b6",
          1224 => x"05",
          1225 => x"a4",
          1226 => x"22",
          1227 => x"08",
          1228 => x"82",
          1229 => x"e4",
          1230 => x"83",
          1231 => x"06",
          1232 => x"72",
          1233 => x"d0",
          1234 => x"a4",
          1235 => x"33",
          1236 => x"70",
          1237 => x"b6",
          1238 => x"05",
          1239 => x"51",
          1240 => x"24",
          1241 => x"b6",
          1242 => x"05",
          1243 => x"06",
          1244 => x"82",
          1245 => x"e4",
          1246 => x"39",
          1247 => x"08",
          1248 => x"53",
          1249 => x"08",
          1250 => x"73",
          1251 => x"54",
          1252 => x"a4",
          1253 => x"34",
          1254 => x"08",
          1255 => x"70",
          1256 => x"81",
          1257 => x"53",
          1258 => x"b1",
          1259 => x"a4",
          1260 => x"33",
          1261 => x"70",
          1262 => x"90",
          1263 => x"2c",
          1264 => x"51",
          1265 => x"82",
          1266 => x"ec",
          1267 => x"75",
          1268 => x"72",
          1269 => x"08",
          1270 => x"af",
          1271 => x"a4",
          1272 => x"33",
          1273 => x"70",
          1274 => x"90",
          1275 => x"2c",
          1276 => x"51",
          1277 => x"82",
          1278 => x"ec",
          1279 => x"75",
          1280 => x"72",
          1281 => x"08",
          1282 => x"82",
          1283 => x"e4",
          1284 => x"83",
          1285 => x"53",
          1286 => x"82",
          1287 => x"ec",
          1288 => x"11",
          1289 => x"82",
          1290 => x"ec",
          1291 => x"90",
          1292 => x"2c",
          1293 => x"73",
          1294 => x"82",
          1295 => x"88",
          1296 => x"a0",
          1297 => x"3f",
          1298 => x"b6",
          1299 => x"05",
          1300 => x"2a",
          1301 => x"51",
          1302 => x"80",
          1303 => x"82",
          1304 => x"88",
          1305 => x"ad",
          1306 => x"3f",
          1307 => x"82",
          1308 => x"e4",
          1309 => x"84",
          1310 => x"06",
          1311 => x"72",
          1312 => x"38",
          1313 => x"08",
          1314 => x"52",
          1315 => x"a5",
          1316 => x"82",
          1317 => x"e4",
          1318 => x"85",
          1319 => x"06",
          1320 => x"72",
          1321 => x"38",
          1322 => x"08",
          1323 => x"52",
          1324 => x"81",
          1325 => x"a4",
          1326 => x"22",
          1327 => x"70",
          1328 => x"51",
          1329 => x"2e",
          1330 => x"b6",
          1331 => x"05",
          1332 => x"51",
          1333 => x"82",
          1334 => x"f4",
          1335 => x"72",
          1336 => x"81",
          1337 => x"82",
          1338 => x"88",
          1339 => x"82",
          1340 => x"f8",
          1341 => x"89",
          1342 => x"b6",
          1343 => x"05",
          1344 => x"2a",
          1345 => x"51",
          1346 => x"80",
          1347 => x"82",
          1348 => x"ec",
          1349 => x"11",
          1350 => x"82",
          1351 => x"ec",
          1352 => x"90",
          1353 => x"2c",
          1354 => x"73",
          1355 => x"82",
          1356 => x"88",
          1357 => x"b0",
          1358 => x"3f",
          1359 => x"b6",
          1360 => x"05",
          1361 => x"2a",
          1362 => x"51",
          1363 => x"80",
          1364 => x"82",
          1365 => x"e8",
          1366 => x"11",
          1367 => x"82",
          1368 => x"e8",
          1369 => x"98",
          1370 => x"2c",
          1371 => x"73",
          1372 => x"82",
          1373 => x"88",
          1374 => x"b0",
          1375 => x"3f",
          1376 => x"b6",
          1377 => x"05",
          1378 => x"2a",
          1379 => x"51",
          1380 => x"b0",
          1381 => x"a4",
          1382 => x"22",
          1383 => x"54",
          1384 => x"a4",
          1385 => x"23",
          1386 => x"70",
          1387 => x"53",
          1388 => x"90",
          1389 => x"a4",
          1390 => x"08",
          1391 => x"87",
          1392 => x"39",
          1393 => x"08",
          1394 => x"53",
          1395 => x"2e",
          1396 => x"97",
          1397 => x"a4",
          1398 => x"08",
          1399 => x"a4",
          1400 => x"33",
          1401 => x"3f",
          1402 => x"82",
          1403 => x"f8",
          1404 => x"72",
          1405 => x"09",
          1406 => x"cb",
          1407 => x"a4",
          1408 => x"22",
          1409 => x"53",
          1410 => x"a4",
          1411 => x"23",
          1412 => x"ff",
          1413 => x"83",
          1414 => x"81",
          1415 => x"b6",
          1416 => x"05",
          1417 => x"b6",
          1418 => x"05",
          1419 => x"52",
          1420 => x"08",
          1421 => x"81",
          1422 => x"a4",
          1423 => x"0c",
          1424 => x"3f",
          1425 => x"82",
          1426 => x"f8",
          1427 => x"72",
          1428 => x"09",
          1429 => x"cb",
          1430 => x"a4",
          1431 => x"22",
          1432 => x"53",
          1433 => x"a4",
          1434 => x"23",
          1435 => x"ff",
          1436 => x"83",
          1437 => x"80",
          1438 => x"b6",
          1439 => x"05",
          1440 => x"b6",
          1441 => x"05",
          1442 => x"52",
          1443 => x"3f",
          1444 => x"08",
          1445 => x"81",
          1446 => x"a4",
          1447 => x"0c",
          1448 => x"82",
          1449 => x"f0",
          1450 => x"b6",
          1451 => x"38",
          1452 => x"08",
          1453 => x"52",
          1454 => x"08",
          1455 => x"ff",
          1456 => x"a4",
          1457 => x"0c",
          1458 => x"08",
          1459 => x"70",
          1460 => x"85",
          1461 => x"39",
          1462 => x"08",
          1463 => x"70",
          1464 => x"81",
          1465 => x"53",
          1466 => x"80",
          1467 => x"b6",
          1468 => x"05",
          1469 => x"54",
          1470 => x"b6",
          1471 => x"05",
          1472 => x"2b",
          1473 => x"51",
          1474 => x"25",
          1475 => x"b6",
          1476 => x"05",
          1477 => x"51",
          1478 => x"d2",
          1479 => x"a4",
          1480 => x"08",
          1481 => x"a4",
          1482 => x"33",
          1483 => x"3f",
          1484 => x"b6",
          1485 => x"05",
          1486 => x"39",
          1487 => x"08",
          1488 => x"53",
          1489 => x"09",
          1490 => x"38",
          1491 => x"b6",
          1492 => x"05",
          1493 => x"82",
          1494 => x"ec",
          1495 => x"0b",
          1496 => x"08",
          1497 => x"8a",
          1498 => x"a4",
          1499 => x"23",
          1500 => x"82",
          1501 => x"88",
          1502 => x"82",
          1503 => x"f8",
          1504 => x"84",
          1505 => x"ea",
          1506 => x"a4",
          1507 => x"08",
          1508 => x"70",
          1509 => x"08",
          1510 => x"51",
          1511 => x"a4",
          1512 => x"08",
          1513 => x"0c",
          1514 => x"82",
          1515 => x"04",
          1516 => x"08",
          1517 => x"a4",
          1518 => x"0d",
          1519 => x"08",
          1520 => x"a4",
          1521 => x"08",
          1522 => x"a4",
          1523 => x"08",
          1524 => x"3f",
          1525 => x"08",
          1526 => x"98",
          1527 => x"3d",
          1528 => x"a4",
          1529 => x"b6",
          1530 => x"82",
          1531 => x"fb",
          1532 => x"0b",
          1533 => x"08",
          1534 => x"82",
          1535 => x"85",
          1536 => x"81",
          1537 => x"32",
          1538 => x"51",
          1539 => x"53",
          1540 => x"8d",
          1541 => x"82",
          1542 => x"f4",
          1543 => x"92",
          1544 => x"a4",
          1545 => x"08",
          1546 => x"82",
          1547 => x"88",
          1548 => x"05",
          1549 => x"08",
          1550 => x"53",
          1551 => x"a4",
          1552 => x"34",
          1553 => x"06",
          1554 => x"2e",
          1555 => x"cd",
          1556 => x"cd",
          1557 => x"82",
          1558 => x"fc",
          1559 => x"90",
          1560 => x"53",
          1561 => x"b6",
          1562 => x"72",
          1563 => x"b1",
          1564 => x"82",
          1565 => x"f8",
          1566 => x"a5",
          1567 => x"ec",
          1568 => x"ec",
          1569 => x"8a",
          1570 => x"08",
          1571 => x"82",
          1572 => x"53",
          1573 => x"8a",
          1574 => x"82",
          1575 => x"f8",
          1576 => x"b6",
          1577 => x"05",
          1578 => x"b6",
          1579 => x"05",
          1580 => x"b6",
          1581 => x"05",
          1582 => x"98",
          1583 => x"0d",
          1584 => x"0c",
          1585 => x"a4",
          1586 => x"b6",
          1587 => x"3d",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"b6",
          1591 => x"05",
          1592 => x"33",
          1593 => x"70",
          1594 => x"81",
          1595 => x"51",
          1596 => x"80",
          1597 => x"ff",
          1598 => x"a4",
          1599 => x"0c",
          1600 => x"82",
          1601 => x"88",
          1602 => x"72",
          1603 => x"a4",
          1604 => x"08",
          1605 => x"b6",
          1606 => x"05",
          1607 => x"82",
          1608 => x"fc",
          1609 => x"81",
          1610 => x"72",
          1611 => x"38",
          1612 => x"08",
          1613 => x"82",
          1614 => x"8c",
          1615 => x"82",
          1616 => x"fc",
          1617 => x"90",
          1618 => x"53",
          1619 => x"b6",
          1620 => x"72",
          1621 => x"ab",
          1622 => x"82",
          1623 => x"f8",
          1624 => x"9f",
          1625 => x"a4",
          1626 => x"08",
          1627 => x"a4",
          1628 => x"0c",
          1629 => x"a4",
          1630 => x"08",
          1631 => x"0c",
          1632 => x"82",
          1633 => x"04",
          1634 => x"08",
          1635 => x"a4",
          1636 => x"0d",
          1637 => x"08",
          1638 => x"a4",
          1639 => x"08",
          1640 => x"82",
          1641 => x"70",
          1642 => x"0c",
          1643 => x"0d",
          1644 => x"0c",
          1645 => x"a4",
          1646 => x"b6",
          1647 => x"3d",
          1648 => x"a4",
          1649 => x"08",
          1650 => x"70",
          1651 => x"81",
          1652 => x"06",
          1653 => x"51",
          1654 => x"2e",
          1655 => x"0b",
          1656 => x"08",
          1657 => x"81",
          1658 => x"b6",
          1659 => x"05",
          1660 => x"33",
          1661 => x"70",
          1662 => x"51",
          1663 => x"80",
          1664 => x"38",
          1665 => x"08",
          1666 => x"82",
          1667 => x"8c",
          1668 => x"54",
          1669 => x"88",
          1670 => x"9f",
          1671 => x"a4",
          1672 => x"08",
          1673 => x"82",
          1674 => x"88",
          1675 => x"57",
          1676 => x"75",
          1677 => x"81",
          1678 => x"82",
          1679 => x"8c",
          1680 => x"11",
          1681 => x"8c",
          1682 => x"b6",
          1683 => x"05",
          1684 => x"b6",
          1685 => x"05",
          1686 => x"80",
          1687 => x"b6",
          1688 => x"05",
          1689 => x"a4",
          1690 => x"08",
          1691 => x"a4",
          1692 => x"08",
          1693 => x"06",
          1694 => x"08",
          1695 => x"72",
          1696 => x"98",
          1697 => x"a3",
          1698 => x"a4",
          1699 => x"08",
          1700 => x"81",
          1701 => x"0c",
          1702 => x"08",
          1703 => x"70",
          1704 => x"08",
          1705 => x"51",
          1706 => x"ff",
          1707 => x"a4",
          1708 => x"0c",
          1709 => x"08",
          1710 => x"82",
          1711 => x"87",
          1712 => x"b6",
          1713 => x"82",
          1714 => x"02",
          1715 => x"0c",
          1716 => x"82",
          1717 => x"88",
          1718 => x"11",
          1719 => x"32",
          1720 => x"51",
          1721 => x"71",
          1722 => x"38",
          1723 => x"b6",
          1724 => x"05",
          1725 => x"39",
          1726 => x"08",
          1727 => x"85",
          1728 => x"86",
          1729 => x"06",
          1730 => x"52",
          1731 => x"80",
          1732 => x"b6",
          1733 => x"05",
          1734 => x"a4",
          1735 => x"08",
          1736 => x"12",
          1737 => x"bf",
          1738 => x"71",
          1739 => x"82",
          1740 => x"88",
          1741 => x"11",
          1742 => x"8c",
          1743 => x"b6",
          1744 => x"05",
          1745 => x"33",
          1746 => x"a4",
          1747 => x"0c",
          1748 => x"82",
          1749 => x"b6",
          1750 => x"05",
          1751 => x"33",
          1752 => x"70",
          1753 => x"51",
          1754 => x"80",
          1755 => x"38",
          1756 => x"08",
          1757 => x"70",
          1758 => x"82",
          1759 => x"fc",
          1760 => x"52",
          1761 => x"08",
          1762 => x"a9",
          1763 => x"a4",
          1764 => x"08",
          1765 => x"08",
          1766 => x"53",
          1767 => x"33",
          1768 => x"51",
          1769 => x"14",
          1770 => x"82",
          1771 => x"f8",
          1772 => x"d7",
          1773 => x"a4",
          1774 => x"08",
          1775 => x"05",
          1776 => x"81",
          1777 => x"b6",
          1778 => x"05",
          1779 => x"a4",
          1780 => x"08",
          1781 => x"08",
          1782 => x"2d",
          1783 => x"08",
          1784 => x"a4",
          1785 => x"0c",
          1786 => x"a4",
          1787 => x"08",
          1788 => x"f2",
          1789 => x"a4",
          1790 => x"08",
          1791 => x"08",
          1792 => x"82",
          1793 => x"88",
          1794 => x"11",
          1795 => x"a4",
          1796 => x"0c",
          1797 => x"a4",
          1798 => x"08",
          1799 => x"81",
          1800 => x"82",
          1801 => x"f0",
          1802 => x"07",
          1803 => x"b6",
          1804 => x"05",
          1805 => x"82",
          1806 => x"f0",
          1807 => x"07",
          1808 => x"b6",
          1809 => x"05",
          1810 => x"a4",
          1811 => x"08",
          1812 => x"a4",
          1813 => x"33",
          1814 => x"ff",
          1815 => x"a4",
          1816 => x"0c",
          1817 => x"b6",
          1818 => x"05",
          1819 => x"08",
          1820 => x"12",
          1821 => x"a4",
          1822 => x"08",
          1823 => x"06",
          1824 => x"a4",
          1825 => x"0c",
          1826 => x"82",
          1827 => x"f8",
          1828 => x"b6",
          1829 => x"3d",
          1830 => x"a4",
          1831 => x"b6",
          1832 => x"82",
          1833 => x"fd",
          1834 => x"b6",
          1835 => x"05",
          1836 => x"a4",
          1837 => x"0c",
          1838 => x"08",
          1839 => x"82",
          1840 => x"f8",
          1841 => x"b6",
          1842 => x"05",
          1843 => x"82",
          1844 => x"b6",
          1845 => x"05",
          1846 => x"a4",
          1847 => x"08",
          1848 => x"38",
          1849 => x"08",
          1850 => x"82",
          1851 => x"90",
          1852 => x"51",
          1853 => x"08",
          1854 => x"71",
          1855 => x"38",
          1856 => x"08",
          1857 => x"82",
          1858 => x"90",
          1859 => x"82",
          1860 => x"fc",
          1861 => x"b6",
          1862 => x"05",
          1863 => x"a4",
          1864 => x"08",
          1865 => x"a4",
          1866 => x"0c",
          1867 => x"08",
          1868 => x"81",
          1869 => x"a4",
          1870 => x"0c",
          1871 => x"08",
          1872 => x"ff",
          1873 => x"a4",
          1874 => x"0c",
          1875 => x"08",
          1876 => x"80",
          1877 => x"38",
          1878 => x"08",
          1879 => x"ff",
          1880 => x"a4",
          1881 => x"0c",
          1882 => x"08",
          1883 => x"ff",
          1884 => x"a4",
          1885 => x"0c",
          1886 => x"08",
          1887 => x"82",
          1888 => x"f8",
          1889 => x"51",
          1890 => x"34",
          1891 => x"82",
          1892 => x"90",
          1893 => x"05",
          1894 => x"08",
          1895 => x"82",
          1896 => x"90",
          1897 => x"05",
          1898 => x"08",
          1899 => x"82",
          1900 => x"90",
          1901 => x"2e",
          1902 => x"b6",
          1903 => x"05",
          1904 => x"33",
          1905 => x"08",
          1906 => x"81",
          1907 => x"a4",
          1908 => x"0c",
          1909 => x"08",
          1910 => x"52",
          1911 => x"34",
          1912 => x"08",
          1913 => x"81",
          1914 => x"a4",
          1915 => x"0c",
          1916 => x"82",
          1917 => x"88",
          1918 => x"82",
          1919 => x"51",
          1920 => x"82",
          1921 => x"04",
          1922 => x"08",
          1923 => x"a4",
          1924 => x"0d",
          1925 => x"08",
          1926 => x"82",
          1927 => x"fc",
          1928 => x"b6",
          1929 => x"05",
          1930 => x"33",
          1931 => x"08",
          1932 => x"81",
          1933 => x"a4",
          1934 => x"0c",
          1935 => x"06",
          1936 => x"80",
          1937 => x"da",
          1938 => x"a4",
          1939 => x"08",
          1940 => x"b6",
          1941 => x"05",
          1942 => x"a4",
          1943 => x"08",
          1944 => x"08",
          1945 => x"31",
          1946 => x"98",
          1947 => x"3d",
          1948 => x"a4",
          1949 => x"b6",
          1950 => x"82",
          1951 => x"fe",
          1952 => x"b6",
          1953 => x"05",
          1954 => x"a4",
          1955 => x"0c",
          1956 => x"08",
          1957 => x"52",
          1958 => x"b6",
          1959 => x"05",
          1960 => x"82",
          1961 => x"8c",
          1962 => x"b6",
          1963 => x"05",
          1964 => x"70",
          1965 => x"b6",
          1966 => x"05",
          1967 => x"82",
          1968 => x"fc",
          1969 => x"81",
          1970 => x"70",
          1971 => x"38",
          1972 => x"82",
          1973 => x"88",
          1974 => x"82",
          1975 => x"51",
          1976 => x"82",
          1977 => x"04",
          1978 => x"08",
          1979 => x"a4",
          1980 => x"0d",
          1981 => x"08",
          1982 => x"82",
          1983 => x"fc",
          1984 => x"b6",
          1985 => x"05",
          1986 => x"a4",
          1987 => x"0c",
          1988 => x"08",
          1989 => x"80",
          1990 => x"38",
          1991 => x"08",
          1992 => x"81",
          1993 => x"a4",
          1994 => x"0c",
          1995 => x"08",
          1996 => x"ff",
          1997 => x"a4",
          1998 => x"0c",
          1999 => x"08",
          2000 => x"80",
          2001 => x"82",
          2002 => x"f8",
          2003 => x"70",
          2004 => x"a4",
          2005 => x"08",
          2006 => x"b6",
          2007 => x"05",
          2008 => x"a4",
          2009 => x"08",
          2010 => x"71",
          2011 => x"a4",
          2012 => x"08",
          2013 => x"b6",
          2014 => x"05",
          2015 => x"39",
          2016 => x"08",
          2017 => x"70",
          2018 => x"0c",
          2019 => x"0d",
          2020 => x"0c",
          2021 => x"a4",
          2022 => x"b6",
          2023 => x"3d",
          2024 => x"a4",
          2025 => x"08",
          2026 => x"f4",
          2027 => x"a4",
          2028 => x"08",
          2029 => x"82",
          2030 => x"8c",
          2031 => x"05",
          2032 => x"08",
          2033 => x"82",
          2034 => x"88",
          2035 => x"33",
          2036 => x"06",
          2037 => x"51",
          2038 => x"84",
          2039 => x"39",
          2040 => x"08",
          2041 => x"52",
          2042 => x"b6",
          2043 => x"05",
          2044 => x"82",
          2045 => x"88",
          2046 => x"81",
          2047 => x"51",
          2048 => x"80",
          2049 => x"a4",
          2050 => x"0c",
          2051 => x"82",
          2052 => x"90",
          2053 => x"05",
          2054 => x"08",
          2055 => x"82",
          2056 => x"90",
          2057 => x"2e",
          2058 => x"81",
          2059 => x"a4",
          2060 => x"08",
          2061 => x"e8",
          2062 => x"a4",
          2063 => x"08",
          2064 => x"53",
          2065 => x"ff",
          2066 => x"a4",
          2067 => x"0c",
          2068 => x"82",
          2069 => x"8c",
          2070 => x"05",
          2071 => x"08",
          2072 => x"82",
          2073 => x"8c",
          2074 => x"33",
          2075 => x"8c",
          2076 => x"82",
          2077 => x"fc",
          2078 => x"39",
          2079 => x"08",
          2080 => x"70",
          2081 => x"a4",
          2082 => x"08",
          2083 => x"71",
          2084 => x"b6",
          2085 => x"05",
          2086 => x"52",
          2087 => x"39",
          2088 => x"b6",
          2089 => x"05",
          2090 => x"a4",
          2091 => x"08",
          2092 => x"0c",
          2093 => x"82",
          2094 => x"04",
          2095 => x"08",
          2096 => x"a4",
          2097 => x"0d",
          2098 => x"08",
          2099 => x"82",
          2100 => x"f8",
          2101 => x"b6",
          2102 => x"05",
          2103 => x"80",
          2104 => x"a4",
          2105 => x"0c",
          2106 => x"82",
          2107 => x"f8",
          2108 => x"71",
          2109 => x"a4",
          2110 => x"08",
          2111 => x"b6",
          2112 => x"05",
          2113 => x"ff",
          2114 => x"70",
          2115 => x"38",
          2116 => x"08",
          2117 => x"ff",
          2118 => x"a4",
          2119 => x"0c",
          2120 => x"08",
          2121 => x"ff",
          2122 => x"ff",
          2123 => x"b6",
          2124 => x"05",
          2125 => x"82",
          2126 => x"f8",
          2127 => x"b6",
          2128 => x"05",
          2129 => x"a4",
          2130 => x"08",
          2131 => x"b6",
          2132 => x"05",
          2133 => x"b6",
          2134 => x"05",
          2135 => x"98",
          2136 => x"0d",
          2137 => x"0c",
          2138 => x"a4",
          2139 => x"b6",
          2140 => x"3d",
          2141 => x"a4",
          2142 => x"08",
          2143 => x"08",
          2144 => x"82",
          2145 => x"90",
          2146 => x"2e",
          2147 => x"82",
          2148 => x"90",
          2149 => x"05",
          2150 => x"08",
          2151 => x"82",
          2152 => x"90",
          2153 => x"05",
          2154 => x"08",
          2155 => x"82",
          2156 => x"90",
          2157 => x"2e",
          2158 => x"b6",
          2159 => x"05",
          2160 => x"82",
          2161 => x"fc",
          2162 => x"52",
          2163 => x"82",
          2164 => x"fc",
          2165 => x"05",
          2166 => x"08",
          2167 => x"ff",
          2168 => x"b6",
          2169 => x"05",
          2170 => x"b6",
          2171 => x"84",
          2172 => x"b6",
          2173 => x"82",
          2174 => x"02",
          2175 => x"0c",
          2176 => x"80",
          2177 => x"a4",
          2178 => x"0c",
          2179 => x"08",
          2180 => x"80",
          2181 => x"82",
          2182 => x"88",
          2183 => x"82",
          2184 => x"88",
          2185 => x"0b",
          2186 => x"08",
          2187 => x"82",
          2188 => x"fc",
          2189 => x"38",
          2190 => x"b6",
          2191 => x"05",
          2192 => x"a4",
          2193 => x"08",
          2194 => x"08",
          2195 => x"82",
          2196 => x"8c",
          2197 => x"25",
          2198 => x"b6",
          2199 => x"05",
          2200 => x"b6",
          2201 => x"05",
          2202 => x"82",
          2203 => x"f0",
          2204 => x"b6",
          2205 => x"05",
          2206 => x"81",
          2207 => x"a4",
          2208 => x"0c",
          2209 => x"08",
          2210 => x"82",
          2211 => x"fc",
          2212 => x"53",
          2213 => x"08",
          2214 => x"52",
          2215 => x"08",
          2216 => x"51",
          2217 => x"82",
          2218 => x"70",
          2219 => x"08",
          2220 => x"54",
          2221 => x"08",
          2222 => x"80",
          2223 => x"82",
          2224 => x"f8",
          2225 => x"82",
          2226 => x"f8",
          2227 => x"b6",
          2228 => x"05",
          2229 => x"b6",
          2230 => x"89",
          2231 => x"b6",
          2232 => x"82",
          2233 => x"02",
          2234 => x"0c",
          2235 => x"80",
          2236 => x"a4",
          2237 => x"0c",
          2238 => x"08",
          2239 => x"80",
          2240 => x"82",
          2241 => x"88",
          2242 => x"82",
          2243 => x"88",
          2244 => x"0b",
          2245 => x"08",
          2246 => x"82",
          2247 => x"8c",
          2248 => x"25",
          2249 => x"b6",
          2250 => x"05",
          2251 => x"b6",
          2252 => x"05",
          2253 => x"82",
          2254 => x"8c",
          2255 => x"82",
          2256 => x"88",
          2257 => x"81",
          2258 => x"b6",
          2259 => x"82",
          2260 => x"f8",
          2261 => x"82",
          2262 => x"fc",
          2263 => x"2e",
          2264 => x"b6",
          2265 => x"05",
          2266 => x"b6",
          2267 => x"05",
          2268 => x"a4",
          2269 => x"08",
          2270 => x"98",
          2271 => x"3d",
          2272 => x"a4",
          2273 => x"b6",
          2274 => x"82",
          2275 => x"fd",
          2276 => x"53",
          2277 => x"08",
          2278 => x"52",
          2279 => x"08",
          2280 => x"51",
          2281 => x"82",
          2282 => x"70",
          2283 => x"0c",
          2284 => x"0d",
          2285 => x"0c",
          2286 => x"a4",
          2287 => x"b6",
          2288 => x"3d",
          2289 => x"82",
          2290 => x"8c",
          2291 => x"82",
          2292 => x"88",
          2293 => x"93",
          2294 => x"98",
          2295 => x"b6",
          2296 => x"85",
          2297 => x"b6",
          2298 => x"82",
          2299 => x"02",
          2300 => x"0c",
          2301 => x"81",
          2302 => x"a4",
          2303 => x"0c",
          2304 => x"b6",
          2305 => x"05",
          2306 => x"a4",
          2307 => x"08",
          2308 => x"08",
          2309 => x"27",
          2310 => x"b6",
          2311 => x"05",
          2312 => x"ae",
          2313 => x"82",
          2314 => x"8c",
          2315 => x"a2",
          2316 => x"a4",
          2317 => x"08",
          2318 => x"a4",
          2319 => x"0c",
          2320 => x"08",
          2321 => x"10",
          2322 => x"08",
          2323 => x"ff",
          2324 => x"b6",
          2325 => x"05",
          2326 => x"80",
          2327 => x"b6",
          2328 => x"05",
          2329 => x"a4",
          2330 => x"08",
          2331 => x"82",
          2332 => x"88",
          2333 => x"b6",
          2334 => x"05",
          2335 => x"b6",
          2336 => x"05",
          2337 => x"a4",
          2338 => x"08",
          2339 => x"08",
          2340 => x"07",
          2341 => x"08",
          2342 => x"82",
          2343 => x"fc",
          2344 => x"2a",
          2345 => x"08",
          2346 => x"82",
          2347 => x"8c",
          2348 => x"2a",
          2349 => x"08",
          2350 => x"ff",
          2351 => x"b6",
          2352 => x"05",
          2353 => x"93",
          2354 => x"a4",
          2355 => x"08",
          2356 => x"a4",
          2357 => x"0c",
          2358 => x"82",
          2359 => x"f8",
          2360 => x"82",
          2361 => x"f4",
          2362 => x"82",
          2363 => x"f4",
          2364 => x"b6",
          2365 => x"3d",
          2366 => x"a4",
          2367 => x"b6",
          2368 => x"82",
          2369 => x"f7",
          2370 => x"0b",
          2371 => x"08",
          2372 => x"82",
          2373 => x"8c",
          2374 => x"80",
          2375 => x"b6",
          2376 => x"05",
          2377 => x"51",
          2378 => x"53",
          2379 => x"a4",
          2380 => x"34",
          2381 => x"06",
          2382 => x"2e",
          2383 => x"91",
          2384 => x"a4",
          2385 => x"08",
          2386 => x"05",
          2387 => x"ce",
          2388 => x"a4",
          2389 => x"33",
          2390 => x"2e",
          2391 => x"a4",
          2392 => x"82",
          2393 => x"f0",
          2394 => x"b6",
          2395 => x"05",
          2396 => x"81",
          2397 => x"70",
          2398 => x"72",
          2399 => x"a4",
          2400 => x"34",
          2401 => x"08",
          2402 => x"53",
          2403 => x"09",
          2404 => x"dc",
          2405 => x"a4",
          2406 => x"08",
          2407 => x"05",
          2408 => x"08",
          2409 => x"33",
          2410 => x"08",
          2411 => x"82",
          2412 => x"f8",
          2413 => x"b6",
          2414 => x"05",
          2415 => x"a4",
          2416 => x"08",
          2417 => x"b6",
          2418 => x"a4",
          2419 => x"08",
          2420 => x"84",
          2421 => x"39",
          2422 => x"b6",
          2423 => x"05",
          2424 => x"a4",
          2425 => x"08",
          2426 => x"05",
          2427 => x"08",
          2428 => x"33",
          2429 => x"08",
          2430 => x"81",
          2431 => x"0b",
          2432 => x"08",
          2433 => x"82",
          2434 => x"88",
          2435 => x"08",
          2436 => x"0c",
          2437 => x"53",
          2438 => x"b6",
          2439 => x"05",
          2440 => x"39",
          2441 => x"08",
          2442 => x"53",
          2443 => x"8d",
          2444 => x"82",
          2445 => x"ec",
          2446 => x"80",
          2447 => x"a4",
          2448 => x"33",
          2449 => x"27",
          2450 => x"b6",
          2451 => x"05",
          2452 => x"b9",
          2453 => x"8d",
          2454 => x"82",
          2455 => x"ec",
          2456 => x"d8",
          2457 => x"82",
          2458 => x"f4",
          2459 => x"39",
          2460 => x"08",
          2461 => x"53",
          2462 => x"90",
          2463 => x"a4",
          2464 => x"33",
          2465 => x"26",
          2466 => x"39",
          2467 => x"b6",
          2468 => x"05",
          2469 => x"39",
          2470 => x"b6",
          2471 => x"05",
          2472 => x"82",
          2473 => x"fc",
          2474 => x"b6",
          2475 => x"05",
          2476 => x"73",
          2477 => x"38",
          2478 => x"08",
          2479 => x"53",
          2480 => x"27",
          2481 => x"b6",
          2482 => x"05",
          2483 => x"51",
          2484 => x"b6",
          2485 => x"05",
          2486 => x"a4",
          2487 => x"33",
          2488 => x"53",
          2489 => x"a4",
          2490 => x"34",
          2491 => x"08",
          2492 => x"53",
          2493 => x"ad",
          2494 => x"a4",
          2495 => x"33",
          2496 => x"53",
          2497 => x"a4",
          2498 => x"34",
          2499 => x"08",
          2500 => x"53",
          2501 => x"8d",
          2502 => x"82",
          2503 => x"ec",
          2504 => x"98",
          2505 => x"a4",
          2506 => x"33",
          2507 => x"08",
          2508 => x"54",
          2509 => x"26",
          2510 => x"0b",
          2511 => x"08",
          2512 => x"80",
          2513 => x"b6",
          2514 => x"05",
          2515 => x"b6",
          2516 => x"05",
          2517 => x"b6",
          2518 => x"05",
          2519 => x"82",
          2520 => x"fc",
          2521 => x"b6",
          2522 => x"05",
          2523 => x"81",
          2524 => x"70",
          2525 => x"52",
          2526 => x"33",
          2527 => x"08",
          2528 => x"fe",
          2529 => x"b6",
          2530 => x"05",
          2531 => x"80",
          2532 => x"82",
          2533 => x"fc",
          2534 => x"82",
          2535 => x"fc",
          2536 => x"b6",
          2537 => x"05",
          2538 => x"a4",
          2539 => x"08",
          2540 => x"81",
          2541 => x"a4",
          2542 => x"0c",
          2543 => x"08",
          2544 => x"82",
          2545 => x"8b",
          2546 => x"b6",
          2547 => x"82",
          2548 => x"02",
          2549 => x"0c",
          2550 => x"80",
          2551 => x"a4",
          2552 => x"34",
          2553 => x"08",
          2554 => x"53",
          2555 => x"82",
          2556 => x"88",
          2557 => x"08",
          2558 => x"33",
          2559 => x"b6",
          2560 => x"05",
          2561 => x"ff",
          2562 => x"a0",
          2563 => x"06",
          2564 => x"b6",
          2565 => x"05",
          2566 => x"81",
          2567 => x"53",
          2568 => x"b6",
          2569 => x"05",
          2570 => x"ad",
          2571 => x"06",
          2572 => x"0b",
          2573 => x"08",
          2574 => x"82",
          2575 => x"88",
          2576 => x"08",
          2577 => x"0c",
          2578 => x"53",
          2579 => x"b6",
          2580 => x"05",
          2581 => x"a4",
          2582 => x"33",
          2583 => x"2e",
          2584 => x"81",
          2585 => x"b6",
          2586 => x"05",
          2587 => x"81",
          2588 => x"70",
          2589 => x"72",
          2590 => x"a4",
          2591 => x"34",
          2592 => x"08",
          2593 => x"82",
          2594 => x"e8",
          2595 => x"b6",
          2596 => x"05",
          2597 => x"2e",
          2598 => x"b6",
          2599 => x"05",
          2600 => x"2e",
          2601 => x"cd",
          2602 => x"82",
          2603 => x"f4",
          2604 => x"b6",
          2605 => x"05",
          2606 => x"81",
          2607 => x"70",
          2608 => x"72",
          2609 => x"a4",
          2610 => x"34",
          2611 => x"82",
          2612 => x"a4",
          2613 => x"34",
          2614 => x"08",
          2615 => x"70",
          2616 => x"71",
          2617 => x"51",
          2618 => x"82",
          2619 => x"f8",
          2620 => x"fe",
          2621 => x"a4",
          2622 => x"33",
          2623 => x"26",
          2624 => x"0b",
          2625 => x"08",
          2626 => x"83",
          2627 => x"b6",
          2628 => x"05",
          2629 => x"73",
          2630 => x"82",
          2631 => x"f8",
          2632 => x"72",
          2633 => x"38",
          2634 => x"0b",
          2635 => x"08",
          2636 => x"82",
          2637 => x"0b",
          2638 => x"08",
          2639 => x"b2",
          2640 => x"a4",
          2641 => x"33",
          2642 => x"27",
          2643 => x"b6",
          2644 => x"05",
          2645 => x"b9",
          2646 => x"8d",
          2647 => x"82",
          2648 => x"ec",
          2649 => x"a5",
          2650 => x"82",
          2651 => x"f4",
          2652 => x"0b",
          2653 => x"08",
          2654 => x"82",
          2655 => x"f8",
          2656 => x"a0",
          2657 => x"cf",
          2658 => x"a4",
          2659 => x"33",
          2660 => x"73",
          2661 => x"82",
          2662 => x"f8",
          2663 => x"11",
          2664 => x"82",
          2665 => x"f8",
          2666 => x"b6",
          2667 => x"05",
          2668 => x"51",
          2669 => x"b6",
          2670 => x"05",
          2671 => x"a4",
          2672 => x"33",
          2673 => x"27",
          2674 => x"b6",
          2675 => x"05",
          2676 => x"51",
          2677 => x"b6",
          2678 => x"05",
          2679 => x"a4",
          2680 => x"33",
          2681 => x"26",
          2682 => x"0b",
          2683 => x"08",
          2684 => x"81",
          2685 => x"b6",
          2686 => x"05",
          2687 => x"a4",
          2688 => x"33",
          2689 => x"74",
          2690 => x"80",
          2691 => x"a4",
          2692 => x"0c",
          2693 => x"82",
          2694 => x"f4",
          2695 => x"82",
          2696 => x"fc",
          2697 => x"82",
          2698 => x"f8",
          2699 => x"12",
          2700 => x"08",
          2701 => x"82",
          2702 => x"88",
          2703 => x"08",
          2704 => x"0c",
          2705 => x"51",
          2706 => x"72",
          2707 => x"a4",
          2708 => x"34",
          2709 => x"82",
          2710 => x"f0",
          2711 => x"72",
          2712 => x"38",
          2713 => x"08",
          2714 => x"30",
          2715 => x"08",
          2716 => x"82",
          2717 => x"8c",
          2718 => x"b6",
          2719 => x"05",
          2720 => x"53",
          2721 => x"b6",
          2722 => x"05",
          2723 => x"a4",
          2724 => x"08",
          2725 => x"0c",
          2726 => x"82",
          2727 => x"04",
          2728 => x"79",
          2729 => x"56",
          2730 => x"80",
          2731 => x"38",
          2732 => x"08",
          2733 => x"3f",
          2734 => x"08",
          2735 => x"85",
          2736 => x"80",
          2737 => x"33",
          2738 => x"2e",
          2739 => x"86",
          2740 => x"55",
          2741 => x"57",
          2742 => x"82",
          2743 => x"70",
          2744 => x"e6",
          2745 => x"b6",
          2746 => x"74",
          2747 => x"51",
          2748 => x"82",
          2749 => x"8b",
          2750 => x"33",
          2751 => x"2e",
          2752 => x"81",
          2753 => x"ff",
          2754 => x"99",
          2755 => x"38",
          2756 => x"82",
          2757 => x"89",
          2758 => x"ff",
          2759 => x"52",
          2760 => x"81",
          2761 => x"84",
          2762 => x"cc",
          2763 => x"08",
          2764 => x"98",
          2765 => x"39",
          2766 => x"51",
          2767 => x"82",
          2768 => x"80",
          2769 => x"9b",
          2770 => x"eb",
          2771 => x"d4",
          2772 => x"39",
          2773 => x"51",
          2774 => x"82",
          2775 => x"80",
          2776 => x"9c",
          2777 => x"cf",
          2778 => x"a0",
          2779 => x"39",
          2780 => x"51",
          2781 => x"82",
          2782 => x"bb",
          2783 => x"ec",
          2784 => x"82",
          2785 => x"af",
          2786 => x"a8",
          2787 => x"82",
          2788 => x"a3",
          2789 => x"d8",
          2790 => x"82",
          2791 => x"97",
          2792 => x"80",
          2793 => x"82",
          2794 => x"8b",
          2795 => x"b0",
          2796 => x"82",
          2797 => x"d8",
          2798 => x"3d",
          2799 => x"3d",
          2800 => x"56",
          2801 => x"e7",
          2802 => x"74",
          2803 => x"e8",
          2804 => x"39",
          2805 => x"74",
          2806 => x"3f",
          2807 => x"08",
          2808 => x"ef",
          2809 => x"b6",
          2810 => x"79",
          2811 => x"82",
          2812 => x"ff",
          2813 => x"87",
          2814 => x"ec",
          2815 => x"02",
          2816 => x"e3",
          2817 => x"57",
          2818 => x"30",
          2819 => x"73",
          2820 => x"59",
          2821 => x"77",
          2822 => x"83",
          2823 => x"74",
          2824 => x"81",
          2825 => x"55",
          2826 => x"81",
          2827 => x"53",
          2828 => x"3d",
          2829 => x"80",
          2830 => x"82",
          2831 => x"57",
          2832 => x"08",
          2833 => x"b6",
          2834 => x"c0",
          2835 => x"82",
          2836 => x"59",
          2837 => x"05",
          2838 => x"53",
          2839 => x"51",
          2840 => x"3f",
          2841 => x"08",
          2842 => x"98",
          2843 => x"7a",
          2844 => x"2e",
          2845 => x"19",
          2846 => x"59",
          2847 => x"3d",
          2848 => x"81",
          2849 => x"76",
          2850 => x"07",
          2851 => x"30",
          2852 => x"72",
          2853 => x"51",
          2854 => x"2e",
          2855 => x"9e",
          2856 => x"c0",
          2857 => x"52",
          2858 => x"92",
          2859 => x"75",
          2860 => x"0c",
          2861 => x"04",
          2862 => x"7d",
          2863 => x"bb",
          2864 => x"5a",
          2865 => x"53",
          2866 => x"51",
          2867 => x"82",
          2868 => x"80",
          2869 => x"80",
          2870 => x"77",
          2871 => x"38",
          2872 => x"cd",
          2873 => x"cd",
          2874 => x"cd",
          2875 => x"cd",
          2876 => x"82",
          2877 => x"53",
          2878 => x"08",
          2879 => x"f8",
          2880 => x"d7",
          2881 => x"e8",
          2882 => x"61",
          2883 => x"98",
          2884 => x"7f",
          2885 => x"82",
          2886 => x"59",
          2887 => x"04",
          2888 => x"98",
          2889 => x"0d",
          2890 => x"0d",
          2891 => x"02",
          2892 => x"cf",
          2893 => x"73",
          2894 => x"5f",
          2895 => x"5e",
          2896 => x"82",
          2897 => x"ff",
          2898 => x"82",
          2899 => x"ff",
          2900 => x"80",
          2901 => x"27",
          2902 => x"7b",
          2903 => x"38",
          2904 => x"a7",
          2905 => x"39",
          2906 => x"72",
          2907 => x"38",
          2908 => x"82",
          2909 => x"ff",
          2910 => x"89",
          2911 => x"c4",
          2912 => x"d7",
          2913 => x"55",
          2914 => x"74",
          2915 => x"7a",
          2916 => x"72",
          2917 => x"9f",
          2918 => x"b8",
          2919 => x"39",
          2920 => x"51",
          2921 => x"3f",
          2922 => x"a1",
          2923 => x"53",
          2924 => x"8e",
          2925 => x"52",
          2926 => x"51",
          2927 => x"3f",
          2928 => x"9f",
          2929 => x"b8",
          2930 => x"15",
          2931 => x"ec",
          2932 => x"51",
          2933 => x"fe",
          2934 => x"9f",
          2935 => x"b7",
          2936 => x"55",
          2937 => x"80",
          2938 => x"18",
          2939 => x"53",
          2940 => x"7a",
          2941 => x"81",
          2942 => x"9f",
          2943 => x"38",
          2944 => x"73",
          2945 => x"ff",
          2946 => x"72",
          2947 => x"38",
          2948 => x"26",
          2949 => x"cd",
          2950 => x"73",
          2951 => x"82",
          2952 => x"52",
          2953 => x"8d",
          2954 => x"55",
          2955 => x"82",
          2956 => x"d3",
          2957 => x"18",
          2958 => x"58",
          2959 => x"82",
          2960 => x"98",
          2961 => x"2c",
          2962 => x"a0",
          2963 => x"06",
          2964 => x"b5",
          2965 => x"98",
          2966 => x"70",
          2967 => x"a0",
          2968 => x"72",
          2969 => x"30",
          2970 => x"73",
          2971 => x"51",
          2972 => x"57",
          2973 => x"73",
          2974 => x"76",
          2975 => x"81",
          2976 => x"80",
          2977 => x"7c",
          2978 => x"78",
          2979 => x"38",
          2980 => x"82",
          2981 => x"8f",
          2982 => x"fc",
          2983 => x"9b",
          2984 => x"9f",
          2985 => x"9f",
          2986 => x"ff",
          2987 => x"82",
          2988 => x"51",
          2989 => x"82",
          2990 => x"82",
          2991 => x"82",
          2992 => x"52",
          2993 => x"51",
          2994 => x"3f",
          2995 => x"84",
          2996 => x"3f",
          2997 => x"04",
          2998 => x"87",
          2999 => x"08",
          3000 => x"3f",
          3001 => x"8e",
          3002 => x"a0",
          3003 => x"3f",
          3004 => x"82",
          3005 => x"2a",
          3006 => x"51",
          3007 => x"2e",
          3008 => x"51",
          3009 => x"82",
          3010 => x"99",
          3011 => x"51",
          3012 => x"72",
          3013 => x"81",
          3014 => x"71",
          3015 => x"38",
          3016 => x"d2",
          3017 => x"c8",
          3018 => x"3f",
          3019 => x"c6",
          3020 => x"2a",
          3021 => x"51",
          3022 => x"2e",
          3023 => x"51",
          3024 => x"82",
          3025 => x"98",
          3026 => x"51",
          3027 => x"72",
          3028 => x"81",
          3029 => x"71",
          3030 => x"38",
          3031 => x"96",
          3032 => x"ec",
          3033 => x"3f",
          3034 => x"8a",
          3035 => x"2a",
          3036 => x"51",
          3037 => x"2e",
          3038 => x"51",
          3039 => x"82",
          3040 => x"98",
          3041 => x"51",
          3042 => x"72",
          3043 => x"81",
          3044 => x"71",
          3045 => x"38",
          3046 => x"da",
          3047 => x"94",
          3048 => x"3f",
          3049 => x"ce",
          3050 => x"2a",
          3051 => x"51",
          3052 => x"2e",
          3053 => x"51",
          3054 => x"82",
          3055 => x"97",
          3056 => x"51",
          3057 => x"72",
          3058 => x"81",
          3059 => x"71",
          3060 => x"38",
          3061 => x"9e",
          3062 => x"bc",
          3063 => x"3f",
          3064 => x"92",
          3065 => x"3f",
          3066 => x"04",
          3067 => x"77",
          3068 => x"a3",
          3069 => x"55",
          3070 => x"52",
          3071 => x"e9",
          3072 => x"82",
          3073 => x"54",
          3074 => x"81",
          3075 => x"f8",
          3076 => x"98",
          3077 => x"89",
          3078 => x"98",
          3079 => x"82",
          3080 => x"07",
          3081 => x"71",
          3082 => x"54",
          3083 => x"82",
          3084 => x"0b",
          3085 => x"94",
          3086 => x"81",
          3087 => x"06",
          3088 => x"cd",
          3089 => x"52",
          3090 => x"b2",
          3091 => x"b6",
          3092 => x"2e",
          3093 => x"b6",
          3094 => x"cf",
          3095 => x"39",
          3096 => x"51",
          3097 => x"3f",
          3098 => x"0b",
          3099 => x"34",
          3100 => x"b1",
          3101 => x"73",
          3102 => x"81",
          3103 => x"82",
          3104 => x"74",
          3105 => x"a9",
          3106 => x"0b",
          3107 => x"0c",
          3108 => x"04",
          3109 => x"80",
          3110 => x"cd",
          3111 => x"5d",
          3112 => x"51",
          3113 => x"3f",
          3114 => x"08",
          3115 => x"59",
          3116 => x"09",
          3117 => x"38",
          3118 => x"83",
          3119 => x"90",
          3120 => x"dc",
          3121 => x"53",
          3122 => x"b7",
          3123 => x"f5",
          3124 => x"b6",
          3125 => x"2e",
          3126 => x"a2",
          3127 => x"a3",
          3128 => x"5f",
          3129 => x"cc",
          3130 => x"ef",
          3131 => x"70",
          3132 => x"f8",
          3133 => x"fd",
          3134 => x"3d",
          3135 => x"51",
          3136 => x"82",
          3137 => x"90",
          3138 => x"2c",
          3139 => x"80",
          3140 => x"a3",
          3141 => x"c2",
          3142 => x"78",
          3143 => x"d2",
          3144 => x"24",
          3145 => x"80",
          3146 => x"38",
          3147 => x"80",
          3148 => x"d4",
          3149 => x"c0",
          3150 => x"38",
          3151 => x"24",
          3152 => x"78",
          3153 => x"8c",
          3154 => x"39",
          3155 => x"2e",
          3156 => x"78",
          3157 => x"92",
          3158 => x"c3",
          3159 => x"38",
          3160 => x"2e",
          3161 => x"8a",
          3162 => x"81",
          3163 => x"86",
          3164 => x"83",
          3165 => x"78",
          3166 => x"89",
          3167 => x"88",
          3168 => x"85",
          3169 => x"38",
          3170 => x"b4",
          3171 => x"11",
          3172 => x"05",
          3173 => x"3f",
          3174 => x"08",
          3175 => x"c5",
          3176 => x"fe",
          3177 => x"ff",
          3178 => x"ec",
          3179 => x"b6",
          3180 => x"2e",
          3181 => x"b4",
          3182 => x"11",
          3183 => x"05",
          3184 => x"3f",
          3185 => x"08",
          3186 => x"b6",
          3187 => x"82",
          3188 => x"ff",
          3189 => x"63",
          3190 => x"79",
          3191 => x"ec",
          3192 => x"78",
          3193 => x"05",
          3194 => x"7a",
          3195 => x"81",
          3196 => x"3d",
          3197 => x"53",
          3198 => x"51",
          3199 => x"82",
          3200 => x"80",
          3201 => x"38",
          3202 => x"fc",
          3203 => x"84",
          3204 => x"bb",
          3205 => x"98",
          3206 => x"fd",
          3207 => x"3d",
          3208 => x"53",
          3209 => x"51",
          3210 => x"82",
          3211 => x"80",
          3212 => x"38",
          3213 => x"51",
          3214 => x"3f",
          3215 => x"63",
          3216 => x"38",
          3217 => x"70",
          3218 => x"33",
          3219 => x"81",
          3220 => x"39",
          3221 => x"80",
          3222 => x"84",
          3223 => x"ef",
          3224 => x"98",
          3225 => x"fc",
          3226 => x"3d",
          3227 => x"53",
          3228 => x"51",
          3229 => x"82",
          3230 => x"80",
          3231 => x"38",
          3232 => x"f8",
          3233 => x"84",
          3234 => x"c3",
          3235 => x"98",
          3236 => x"fc",
          3237 => x"a2",
          3238 => x"ae",
          3239 => x"5a",
          3240 => x"a8",
          3241 => x"33",
          3242 => x"5a",
          3243 => x"2e",
          3244 => x"55",
          3245 => x"33",
          3246 => x"82",
          3247 => x"ff",
          3248 => x"81",
          3249 => x"05",
          3250 => x"39",
          3251 => x"b8",
          3252 => x"39",
          3253 => x"80",
          3254 => x"84",
          3255 => x"ef",
          3256 => x"98",
          3257 => x"38",
          3258 => x"33",
          3259 => x"2e",
          3260 => x"b4",
          3261 => x"80",
          3262 => x"b5",
          3263 => x"78",
          3264 => x"38",
          3265 => x"08",
          3266 => x"82",
          3267 => x"59",
          3268 => x"88",
          3269 => x"cc",
          3270 => x"39",
          3271 => x"33",
          3272 => x"2e",
          3273 => x"b4",
          3274 => x"9a",
          3275 => x"82",
          3276 => x"80",
          3277 => x"82",
          3278 => x"44",
          3279 => x"b4",
          3280 => x"80",
          3281 => x"3d",
          3282 => x"53",
          3283 => x"51",
          3284 => x"82",
          3285 => x"80",
          3286 => x"b5",
          3287 => x"78",
          3288 => x"38",
          3289 => x"08",
          3290 => x"39",
          3291 => x"33",
          3292 => x"2e",
          3293 => x"b4",
          3294 => x"bb",
          3295 => x"86",
          3296 => x"80",
          3297 => x"82",
          3298 => x"43",
          3299 => x"b5",
          3300 => x"78",
          3301 => x"38",
          3302 => x"08",
          3303 => x"82",
          3304 => x"59",
          3305 => x"88",
          3306 => x"e0",
          3307 => x"39",
          3308 => x"08",
          3309 => x"b4",
          3310 => x"11",
          3311 => x"05",
          3312 => x"3f",
          3313 => x"08",
          3314 => x"38",
          3315 => x"5c",
          3316 => x"83",
          3317 => x"7a",
          3318 => x"30",
          3319 => x"9f",
          3320 => x"06",
          3321 => x"5a",
          3322 => x"88",
          3323 => x"2e",
          3324 => x"42",
          3325 => x"51",
          3326 => x"a0",
          3327 => x"61",
          3328 => x"63",
          3329 => x"3f",
          3330 => x"51",
          3331 => x"b4",
          3332 => x"11",
          3333 => x"05",
          3334 => x"3f",
          3335 => x"08",
          3336 => x"c1",
          3337 => x"fe",
          3338 => x"ff",
          3339 => x"e7",
          3340 => x"b6",
          3341 => x"2e",
          3342 => x"59",
          3343 => x"05",
          3344 => x"63",
          3345 => x"b4",
          3346 => x"11",
          3347 => x"05",
          3348 => x"3f",
          3349 => x"08",
          3350 => x"89",
          3351 => x"33",
          3352 => x"a3",
          3353 => x"aa",
          3354 => x"cd",
          3355 => x"80",
          3356 => x"51",
          3357 => x"3f",
          3358 => x"33",
          3359 => x"2e",
          3360 => x"9f",
          3361 => x"38",
          3362 => x"fc",
          3363 => x"84",
          3364 => x"bb",
          3365 => x"98",
          3366 => x"91",
          3367 => x"02",
          3368 => x"33",
          3369 => x"81",
          3370 => x"b1",
          3371 => x"bc",
          3372 => x"3f",
          3373 => x"b4",
          3374 => x"11",
          3375 => x"05",
          3376 => x"3f",
          3377 => x"08",
          3378 => x"99",
          3379 => x"fe",
          3380 => x"ff",
          3381 => x"e0",
          3382 => x"b6",
          3383 => x"2e",
          3384 => x"59",
          3385 => x"22",
          3386 => x"05",
          3387 => x"41",
          3388 => x"f0",
          3389 => x"84",
          3390 => x"82",
          3391 => x"98",
          3392 => x"f7",
          3393 => x"70",
          3394 => x"82",
          3395 => x"ff",
          3396 => x"82",
          3397 => x"53",
          3398 => x"79",
          3399 => x"90",
          3400 => x"79",
          3401 => x"ae",
          3402 => x"38",
          3403 => x"87",
          3404 => x"05",
          3405 => x"b4",
          3406 => x"11",
          3407 => x"05",
          3408 => x"3f",
          3409 => x"08",
          3410 => x"38",
          3411 => x"be",
          3412 => x"70",
          3413 => x"23",
          3414 => x"aa",
          3415 => x"bc",
          3416 => x"3f",
          3417 => x"b4",
          3418 => x"11",
          3419 => x"05",
          3420 => x"3f",
          3421 => x"08",
          3422 => x"e9",
          3423 => x"fe",
          3424 => x"ff",
          3425 => x"de",
          3426 => x"b6",
          3427 => x"2e",
          3428 => x"60",
          3429 => x"60",
          3430 => x"b4",
          3431 => x"11",
          3432 => x"05",
          3433 => x"3f",
          3434 => x"08",
          3435 => x"b5",
          3436 => x"08",
          3437 => x"a3",
          3438 => x"a8",
          3439 => x"cd",
          3440 => x"80",
          3441 => x"51",
          3442 => x"3f",
          3443 => x"33",
          3444 => x"2e",
          3445 => x"9f",
          3446 => x"38",
          3447 => x"f0",
          3448 => x"84",
          3449 => x"96",
          3450 => x"98",
          3451 => x"8d",
          3452 => x"71",
          3453 => x"84",
          3454 => x"b5",
          3455 => x"bc",
          3456 => x"3f",
          3457 => x"b4",
          3458 => x"11",
          3459 => x"05",
          3460 => x"3f",
          3461 => x"08",
          3462 => x"c9",
          3463 => x"82",
          3464 => x"ff",
          3465 => x"63",
          3466 => x"b4",
          3467 => x"11",
          3468 => x"05",
          3469 => x"3f",
          3470 => x"08",
          3471 => x"a5",
          3472 => x"82",
          3473 => x"ff",
          3474 => x"63",
          3475 => x"82",
          3476 => x"80",
          3477 => x"38",
          3478 => x"08",
          3479 => x"94",
          3480 => x"f7",
          3481 => x"39",
          3482 => x"51",
          3483 => x"ff",
          3484 => x"f4",
          3485 => x"a4",
          3486 => x"ea",
          3487 => x"ff",
          3488 => x"a7",
          3489 => x"39",
          3490 => x"33",
          3491 => x"2e",
          3492 => x"7d",
          3493 => x"78",
          3494 => x"cf",
          3495 => x"ff",
          3496 => x"83",
          3497 => x"b6",
          3498 => x"81",
          3499 => x"2e",
          3500 => x"82",
          3501 => x"7a",
          3502 => x"38",
          3503 => x"7a",
          3504 => x"38",
          3505 => x"82",
          3506 => x"7b",
          3507 => x"e4",
          3508 => x"82",
          3509 => x"b4",
          3510 => x"05",
          3511 => x"e3",
          3512 => x"7b",
          3513 => x"ff",
          3514 => x"cf",
          3515 => x"39",
          3516 => x"a4",
          3517 => x"53",
          3518 => x"52",
          3519 => x"b0",
          3520 => x"a8",
          3521 => x"39",
          3522 => x"53",
          3523 => x"52",
          3524 => x"b0",
          3525 => x"a8",
          3526 => x"b4",
          3527 => x"b6",
          3528 => x"56",
          3529 => x"54",
          3530 => x"53",
          3531 => x"52",
          3532 => x"b0",
          3533 => x"80",
          3534 => x"98",
          3535 => x"98",
          3536 => x"30",
          3537 => x"80",
          3538 => x"5b",
          3539 => x"7a",
          3540 => x"38",
          3541 => x"7a",
          3542 => x"80",
          3543 => x"81",
          3544 => x"ff",
          3545 => x"7a",
          3546 => x"7d",
          3547 => x"81",
          3548 => x"78",
          3549 => x"ff",
          3550 => x"06",
          3551 => x"82",
          3552 => x"c0",
          3553 => x"dd",
          3554 => x"0d",
          3555 => x"b6",
          3556 => x"c0",
          3557 => x"08",
          3558 => x"84",
          3559 => x"51",
          3560 => x"82",
          3561 => x"90",
          3562 => x"55",
          3563 => x"80",
          3564 => x"d7",
          3565 => x"82",
          3566 => x"07",
          3567 => x"c0",
          3568 => x"08",
          3569 => x"84",
          3570 => x"51",
          3571 => x"82",
          3572 => x"90",
          3573 => x"55",
          3574 => x"80",
          3575 => x"d7",
          3576 => x"82",
          3577 => x"07",
          3578 => x"80",
          3579 => x"c0",
          3580 => x"8c",
          3581 => x"87",
          3582 => x"0c",
          3583 => x"5a",
          3584 => x"5b",
          3585 => x"05",
          3586 => x"80",
          3587 => x"e8",
          3588 => x"70",
          3589 => x"70",
          3590 => x"cd",
          3591 => x"89",
          3592 => x"ff",
          3593 => x"9c",
          3594 => x"ba",
          3595 => x"a8",
          3596 => x"b2",
          3597 => x"d5",
          3598 => x"3f",
          3599 => x"db",
          3600 => x"3f",
          3601 => x"3d",
          3602 => x"83",
          3603 => x"2b",
          3604 => x"3f",
          3605 => x"08",
          3606 => x"72",
          3607 => x"54",
          3608 => x"25",
          3609 => x"82",
          3610 => x"84",
          3611 => x"fc",
          3612 => x"70",
          3613 => x"80",
          3614 => x"72",
          3615 => x"8a",
          3616 => x"51",
          3617 => x"09",
          3618 => x"38",
          3619 => x"f1",
          3620 => x"51",
          3621 => x"09",
          3622 => x"38",
          3623 => x"81",
          3624 => x"73",
          3625 => x"81",
          3626 => x"84",
          3627 => x"52",
          3628 => x"52",
          3629 => x"2e",
          3630 => x"54",
          3631 => x"9d",
          3632 => x"38",
          3633 => x"12",
          3634 => x"33",
          3635 => x"a0",
          3636 => x"81",
          3637 => x"2e",
          3638 => x"ea",
          3639 => x"33",
          3640 => x"a0",
          3641 => x"06",
          3642 => x"54",
          3643 => x"70",
          3644 => x"25",
          3645 => x"51",
          3646 => x"2e",
          3647 => x"72",
          3648 => x"54",
          3649 => x"0c",
          3650 => x"82",
          3651 => x"86",
          3652 => x"fc",
          3653 => x"53",
          3654 => x"2e",
          3655 => x"3d",
          3656 => x"72",
          3657 => x"3f",
          3658 => x"08",
          3659 => x"53",
          3660 => x"53",
          3661 => x"98",
          3662 => x"0d",
          3663 => x"0d",
          3664 => x"33",
          3665 => x"53",
          3666 => x"8b",
          3667 => x"38",
          3668 => x"ff",
          3669 => x"52",
          3670 => x"81",
          3671 => x"13",
          3672 => x"52",
          3673 => x"80",
          3674 => x"13",
          3675 => x"52",
          3676 => x"80",
          3677 => x"13",
          3678 => x"52",
          3679 => x"80",
          3680 => x"13",
          3681 => x"52",
          3682 => x"26",
          3683 => x"8a",
          3684 => x"87",
          3685 => x"e7",
          3686 => x"38",
          3687 => x"c0",
          3688 => x"72",
          3689 => x"98",
          3690 => x"13",
          3691 => x"98",
          3692 => x"13",
          3693 => x"98",
          3694 => x"13",
          3695 => x"98",
          3696 => x"13",
          3697 => x"98",
          3698 => x"13",
          3699 => x"98",
          3700 => x"87",
          3701 => x"0c",
          3702 => x"98",
          3703 => x"0b",
          3704 => x"9c",
          3705 => x"71",
          3706 => x"0c",
          3707 => x"04",
          3708 => x"7f",
          3709 => x"98",
          3710 => x"7d",
          3711 => x"98",
          3712 => x"7d",
          3713 => x"c0",
          3714 => x"5a",
          3715 => x"34",
          3716 => x"b4",
          3717 => x"83",
          3718 => x"c0",
          3719 => x"5a",
          3720 => x"34",
          3721 => x"ac",
          3722 => x"85",
          3723 => x"c0",
          3724 => x"5a",
          3725 => x"34",
          3726 => x"a4",
          3727 => x"88",
          3728 => x"c0",
          3729 => x"5a",
          3730 => x"23",
          3731 => x"79",
          3732 => x"06",
          3733 => x"ff",
          3734 => x"86",
          3735 => x"85",
          3736 => x"84",
          3737 => x"83",
          3738 => x"82",
          3739 => x"7d",
          3740 => x"06",
          3741 => x"c0",
          3742 => x"df",
          3743 => x"0d",
          3744 => x"0d",
          3745 => x"33",
          3746 => x"33",
          3747 => x"06",
          3748 => x"87",
          3749 => x"51",
          3750 => x"86",
          3751 => x"94",
          3752 => x"08",
          3753 => x"70",
          3754 => x"54",
          3755 => x"2e",
          3756 => x"91",
          3757 => x"06",
          3758 => x"d7",
          3759 => x"32",
          3760 => x"51",
          3761 => x"2e",
          3762 => x"93",
          3763 => x"06",
          3764 => x"ff",
          3765 => x"81",
          3766 => x"87",
          3767 => x"52",
          3768 => x"86",
          3769 => x"94",
          3770 => x"72",
          3771 => x"b6",
          3772 => x"3d",
          3773 => x"3d",
          3774 => x"05",
          3775 => x"70",
          3776 => x"52",
          3777 => x"b4",
          3778 => x"3d",
          3779 => x"3d",
          3780 => x"05",
          3781 => x"8a",
          3782 => x"06",
          3783 => x"52",
          3784 => x"3f",
          3785 => x"33",
          3786 => x"06",
          3787 => x"c0",
          3788 => x"76",
          3789 => x"38",
          3790 => x"94",
          3791 => x"70",
          3792 => x"81",
          3793 => x"54",
          3794 => x"8c",
          3795 => x"2a",
          3796 => x"51",
          3797 => x"38",
          3798 => x"70",
          3799 => x"53",
          3800 => x"8d",
          3801 => x"2a",
          3802 => x"51",
          3803 => x"be",
          3804 => x"ff",
          3805 => x"c0",
          3806 => x"72",
          3807 => x"38",
          3808 => x"90",
          3809 => x"0c",
          3810 => x"b6",
          3811 => x"3d",
          3812 => x"3d",
          3813 => x"80",
          3814 => x"81",
          3815 => x"53",
          3816 => x"2e",
          3817 => x"71",
          3818 => x"81",
          3819 => x"b8",
          3820 => x"ff",
          3821 => x"55",
          3822 => x"94",
          3823 => x"80",
          3824 => x"87",
          3825 => x"51",
          3826 => x"96",
          3827 => x"06",
          3828 => x"70",
          3829 => x"38",
          3830 => x"70",
          3831 => x"51",
          3832 => x"72",
          3833 => x"81",
          3834 => x"70",
          3835 => x"38",
          3836 => x"70",
          3837 => x"51",
          3838 => x"38",
          3839 => x"06",
          3840 => x"94",
          3841 => x"80",
          3842 => x"87",
          3843 => x"52",
          3844 => x"81",
          3845 => x"70",
          3846 => x"53",
          3847 => x"ff",
          3848 => x"82",
          3849 => x"89",
          3850 => x"fe",
          3851 => x"b4",
          3852 => x"81",
          3853 => x"52",
          3854 => x"84",
          3855 => x"2e",
          3856 => x"c0",
          3857 => x"70",
          3858 => x"2a",
          3859 => x"51",
          3860 => x"80",
          3861 => x"71",
          3862 => x"51",
          3863 => x"80",
          3864 => x"2e",
          3865 => x"c0",
          3866 => x"71",
          3867 => x"ff",
          3868 => x"98",
          3869 => x"3d",
          3870 => x"af",
          3871 => x"98",
          3872 => x"06",
          3873 => x"0c",
          3874 => x"0d",
          3875 => x"33",
          3876 => x"06",
          3877 => x"c0",
          3878 => x"70",
          3879 => x"38",
          3880 => x"94",
          3881 => x"70",
          3882 => x"81",
          3883 => x"51",
          3884 => x"80",
          3885 => x"72",
          3886 => x"51",
          3887 => x"80",
          3888 => x"2e",
          3889 => x"c0",
          3890 => x"71",
          3891 => x"2b",
          3892 => x"51",
          3893 => x"82",
          3894 => x"84",
          3895 => x"ff",
          3896 => x"c0",
          3897 => x"70",
          3898 => x"06",
          3899 => x"80",
          3900 => x"38",
          3901 => x"a4",
          3902 => x"bc",
          3903 => x"9e",
          3904 => x"b4",
          3905 => x"c0",
          3906 => x"82",
          3907 => x"87",
          3908 => x"08",
          3909 => x"0c",
          3910 => x"9c",
          3911 => x"cc",
          3912 => x"9e",
          3913 => x"b4",
          3914 => x"c0",
          3915 => x"82",
          3916 => x"87",
          3917 => x"08",
          3918 => x"0c",
          3919 => x"b4",
          3920 => x"dc",
          3921 => x"9e",
          3922 => x"b4",
          3923 => x"c0",
          3924 => x"82",
          3925 => x"87",
          3926 => x"08",
          3927 => x"0c",
          3928 => x"c4",
          3929 => x"ec",
          3930 => x"9e",
          3931 => x"70",
          3932 => x"23",
          3933 => x"84",
          3934 => x"f4",
          3935 => x"9e",
          3936 => x"b4",
          3937 => x"c0",
          3938 => x"82",
          3939 => x"81",
          3940 => x"80",
          3941 => x"87",
          3942 => x"08",
          3943 => x"0a",
          3944 => x"52",
          3945 => x"83",
          3946 => x"71",
          3947 => x"34",
          3948 => x"c0",
          3949 => x"70",
          3950 => x"06",
          3951 => x"70",
          3952 => x"38",
          3953 => x"82",
          3954 => x"80",
          3955 => x"9e",
          3956 => x"90",
          3957 => x"51",
          3958 => x"80",
          3959 => x"81",
          3960 => x"b5",
          3961 => x"0b",
          3962 => x"90",
          3963 => x"80",
          3964 => x"52",
          3965 => x"2e",
          3966 => x"52",
          3967 => x"84",
          3968 => x"87",
          3969 => x"08",
          3970 => x"80",
          3971 => x"52",
          3972 => x"83",
          3973 => x"71",
          3974 => x"34",
          3975 => x"c0",
          3976 => x"70",
          3977 => x"06",
          3978 => x"70",
          3979 => x"38",
          3980 => x"82",
          3981 => x"80",
          3982 => x"9e",
          3983 => x"84",
          3984 => x"51",
          3985 => x"80",
          3986 => x"81",
          3987 => x"b5",
          3988 => x"0b",
          3989 => x"90",
          3990 => x"80",
          3991 => x"52",
          3992 => x"2e",
          3993 => x"52",
          3994 => x"88",
          3995 => x"87",
          3996 => x"08",
          3997 => x"80",
          3998 => x"52",
          3999 => x"83",
          4000 => x"71",
          4001 => x"34",
          4002 => x"c0",
          4003 => x"70",
          4004 => x"06",
          4005 => x"70",
          4006 => x"38",
          4007 => x"82",
          4008 => x"80",
          4009 => x"9e",
          4010 => x"a0",
          4011 => x"52",
          4012 => x"2e",
          4013 => x"52",
          4014 => x"8b",
          4015 => x"9e",
          4016 => x"98",
          4017 => x"8a",
          4018 => x"51",
          4019 => x"8c",
          4020 => x"87",
          4021 => x"08",
          4022 => x"06",
          4023 => x"70",
          4024 => x"38",
          4025 => x"82",
          4026 => x"87",
          4027 => x"08",
          4028 => x"06",
          4029 => x"51",
          4030 => x"82",
          4031 => x"80",
          4032 => x"9e",
          4033 => x"88",
          4034 => x"52",
          4035 => x"83",
          4036 => x"71",
          4037 => x"34",
          4038 => x"90",
          4039 => x"06",
          4040 => x"82",
          4041 => x"83",
          4042 => x"fb",
          4043 => x"a5",
          4044 => x"95",
          4045 => x"b5",
          4046 => x"73",
          4047 => x"38",
          4048 => x"51",
          4049 => x"3f",
          4050 => x"51",
          4051 => x"3f",
          4052 => x"33",
          4053 => x"2e",
          4054 => x"b4",
          4055 => x"b4",
          4056 => x"54",
          4057 => x"98",
          4058 => x"ef",
          4059 => x"87",
          4060 => x"80",
          4061 => x"82",
          4062 => x"82",
          4063 => x"11",
          4064 => x"a6",
          4065 => x"94",
          4066 => x"b5",
          4067 => x"73",
          4068 => x"38",
          4069 => x"08",
          4070 => x"08",
          4071 => x"82",
          4072 => x"ff",
          4073 => x"82",
          4074 => x"54",
          4075 => x"94",
          4076 => x"c4",
          4077 => x"c8",
          4078 => x"52",
          4079 => x"51",
          4080 => x"3f",
          4081 => x"33",
          4082 => x"2e",
          4083 => x"b4",
          4084 => x"b4",
          4085 => x"54",
          4086 => x"88",
          4087 => x"fb",
          4088 => x"8b",
          4089 => x"80",
          4090 => x"82",
          4091 => x"52",
          4092 => x"51",
          4093 => x"3f",
          4094 => x"33",
          4095 => x"2e",
          4096 => x"b5",
          4097 => x"82",
          4098 => x"ff",
          4099 => x"82",
          4100 => x"54",
          4101 => x"8e",
          4102 => x"8e",
          4103 => x"a7",
          4104 => x"93",
          4105 => x"b5",
          4106 => x"73",
          4107 => x"38",
          4108 => x"51",
          4109 => x"3f",
          4110 => x"33",
          4111 => x"2e",
          4112 => x"a8",
          4113 => x"af",
          4114 => x"b5",
          4115 => x"73",
          4116 => x"38",
          4117 => x"51",
          4118 => x"3f",
          4119 => x"33",
          4120 => x"2e",
          4121 => x"a8",
          4122 => x"ae",
          4123 => x"b5",
          4124 => x"73",
          4125 => x"38",
          4126 => x"51",
          4127 => x"3f",
          4128 => x"51",
          4129 => x"3f",
          4130 => x"08",
          4131 => x"cc",
          4132 => x"c7",
          4133 => x"e8",
          4134 => x"a8",
          4135 => x"92",
          4136 => x"b4",
          4137 => x"82",
          4138 => x"ff",
          4139 => x"82",
          4140 => x"ff",
          4141 => x"82",
          4142 => x"52",
          4143 => x"51",
          4144 => x"3f",
          4145 => x"08",
          4146 => x"c0",
          4147 => x"c5",
          4148 => x"b6",
          4149 => x"84",
          4150 => x"71",
          4151 => x"82",
          4152 => x"52",
          4153 => x"51",
          4154 => x"3f",
          4155 => x"33",
          4156 => x"2e",
          4157 => x"b4",
          4158 => x"bd",
          4159 => x"75",
          4160 => x"3f",
          4161 => x"08",
          4162 => x"29",
          4163 => x"54",
          4164 => x"98",
          4165 => x"aa",
          4166 => x"91",
          4167 => x"b5",
          4168 => x"73",
          4169 => x"38",
          4170 => x"08",
          4171 => x"c0",
          4172 => x"c4",
          4173 => x"b6",
          4174 => x"84",
          4175 => x"71",
          4176 => x"82",
          4177 => x"52",
          4178 => x"51",
          4179 => x"3f",
          4180 => x"b0",
          4181 => x"3d",
          4182 => x"3d",
          4183 => x"05",
          4184 => x"52",
          4185 => x"aa",
          4186 => x"29",
          4187 => x"05",
          4188 => x"04",
          4189 => x"51",
          4190 => x"ab",
          4191 => x"39",
          4192 => x"51",
          4193 => x"ab",
          4194 => x"39",
          4195 => x"51",
          4196 => x"ab",
          4197 => x"90",
          4198 => x"3d",
          4199 => x"88",
          4200 => x"80",
          4201 => x"96",
          4202 => x"82",
          4203 => x"87",
          4204 => x"0c",
          4205 => x"0d",
          4206 => x"70",
          4207 => x"98",
          4208 => x"2c",
          4209 => x"70",
          4210 => x"53",
          4211 => x"51",
          4212 => x"ab",
          4213 => x"55",
          4214 => x"25",
          4215 => x"ab",
          4216 => x"12",
          4217 => x"97",
          4218 => x"33",
          4219 => x"70",
          4220 => x"81",
          4221 => x"81",
          4222 => x"b6",
          4223 => x"3d",
          4224 => x"3d",
          4225 => x"84",
          4226 => x"33",
          4227 => x"56",
          4228 => x"2e",
          4229 => x"cd",
          4230 => x"88",
          4231 => x"95",
          4232 => x"ec",
          4233 => x"51",
          4234 => x"3f",
          4235 => x"08",
          4236 => x"ff",
          4237 => x"73",
          4238 => x"53",
          4239 => x"72",
          4240 => x"53",
          4241 => x"51",
          4242 => x"3f",
          4243 => x"87",
          4244 => x"f6",
          4245 => x"02",
          4246 => x"05",
          4247 => x"05",
          4248 => x"82",
          4249 => x"70",
          4250 => x"b5",
          4251 => x"08",
          4252 => x"5a",
          4253 => x"80",
          4254 => x"74",
          4255 => x"3f",
          4256 => x"33",
          4257 => x"82",
          4258 => x"81",
          4259 => x"58",
          4260 => x"fb",
          4261 => x"98",
          4262 => x"82",
          4263 => x"70",
          4264 => x"b5",
          4265 => x"08",
          4266 => x"74",
          4267 => x"38",
          4268 => x"52",
          4269 => x"b8",
          4270 => x"b5",
          4271 => x"05",
          4272 => x"b5",
          4273 => x"81",
          4274 => x"93",
          4275 => x"38",
          4276 => x"b5",
          4277 => x"80",
          4278 => x"82",
          4279 => x"56",
          4280 => x"ac",
          4281 => x"e8",
          4282 => x"a4",
          4283 => x"fc",
          4284 => x"53",
          4285 => x"51",
          4286 => x"3f",
          4287 => x"08",
          4288 => x"81",
          4289 => x"82",
          4290 => x"51",
          4291 => x"3f",
          4292 => x"04",
          4293 => x"82",
          4294 => x"93",
          4295 => x"52",
          4296 => x"89",
          4297 => x"99",
          4298 => x"73",
          4299 => x"84",
          4300 => x"73",
          4301 => x"38",
          4302 => x"b5",
          4303 => x"b5",
          4304 => x"71",
          4305 => x"38",
          4306 => x"de",
          4307 => x"b5",
          4308 => x"99",
          4309 => x"0b",
          4310 => x"0c",
          4311 => x"04",
          4312 => x"81",
          4313 => x"82",
          4314 => x"51",
          4315 => x"3f",
          4316 => x"08",
          4317 => x"82",
          4318 => x"53",
          4319 => x"88",
          4320 => x"56",
          4321 => x"3f",
          4322 => x"08",
          4323 => x"38",
          4324 => x"b4",
          4325 => x"b6",
          4326 => x"80",
          4327 => x"98",
          4328 => x"38",
          4329 => x"08",
          4330 => x"17",
          4331 => x"74",
          4332 => x"76",
          4333 => x"82",
          4334 => x"57",
          4335 => x"3f",
          4336 => x"09",
          4337 => x"af",
          4338 => x"0d",
          4339 => x"0d",
          4340 => x"ad",
          4341 => x"5a",
          4342 => x"58",
          4343 => x"b5",
          4344 => x"80",
          4345 => x"82",
          4346 => x"81",
          4347 => x"0b",
          4348 => x"08",
          4349 => x"f8",
          4350 => x"70",
          4351 => x"8b",
          4352 => x"b6",
          4353 => x"2e",
          4354 => x"51",
          4355 => x"3f",
          4356 => x"08",
          4357 => x"55",
          4358 => x"b6",
          4359 => x"8e",
          4360 => x"98",
          4361 => x"70",
          4362 => x"80",
          4363 => x"09",
          4364 => x"72",
          4365 => x"51",
          4366 => x"77",
          4367 => x"73",
          4368 => x"82",
          4369 => x"8c",
          4370 => x"51",
          4371 => x"3f",
          4372 => x"08",
          4373 => x"38",
          4374 => x"51",
          4375 => x"3f",
          4376 => x"09",
          4377 => x"38",
          4378 => x"51",
          4379 => x"3f",
          4380 => x"b3",
          4381 => x"3d",
          4382 => x"b6",
          4383 => x"34",
          4384 => x"82",
          4385 => x"a9",
          4386 => x"f6",
          4387 => x"7e",
          4388 => x"72",
          4389 => x"5a",
          4390 => x"2e",
          4391 => x"a2",
          4392 => x"78",
          4393 => x"76",
          4394 => x"81",
          4395 => x"70",
          4396 => x"58",
          4397 => x"2e",
          4398 => x"86",
          4399 => x"26",
          4400 => x"54",
          4401 => x"82",
          4402 => x"70",
          4403 => x"ff",
          4404 => x"82",
          4405 => x"53",
          4406 => x"08",
          4407 => x"b5",
          4408 => x"98",
          4409 => x"38",
          4410 => x"55",
          4411 => x"88",
          4412 => x"2e",
          4413 => x"39",
          4414 => x"ac",
          4415 => x"5a",
          4416 => x"11",
          4417 => x"51",
          4418 => x"82",
          4419 => x"80",
          4420 => x"ff",
          4421 => x"52",
          4422 => x"b1",
          4423 => x"98",
          4424 => x"06",
          4425 => x"38",
          4426 => x"39",
          4427 => x"81",
          4428 => x"54",
          4429 => x"ff",
          4430 => x"54",
          4431 => x"98",
          4432 => x"0d",
          4433 => x"0d",
          4434 => x"b2",
          4435 => x"3d",
          4436 => x"5a",
          4437 => x"3d",
          4438 => x"f0",
          4439 => x"ec",
          4440 => x"73",
          4441 => x"73",
          4442 => x"33",
          4443 => x"83",
          4444 => x"76",
          4445 => x"bc",
          4446 => x"76",
          4447 => x"73",
          4448 => x"ad",
          4449 => x"98",
          4450 => x"b6",
          4451 => x"b5",
          4452 => x"b6",
          4453 => x"2e",
          4454 => x"93",
          4455 => x"82",
          4456 => x"51",
          4457 => x"3f",
          4458 => x"08",
          4459 => x"38",
          4460 => x"51",
          4461 => x"3f",
          4462 => x"82",
          4463 => x"5b",
          4464 => x"08",
          4465 => x"52",
          4466 => x"52",
          4467 => x"b7",
          4468 => x"98",
          4469 => x"b6",
          4470 => x"2e",
          4471 => x"80",
          4472 => x"b6",
          4473 => x"ff",
          4474 => x"82",
          4475 => x"55",
          4476 => x"b6",
          4477 => x"a9",
          4478 => x"98",
          4479 => x"70",
          4480 => x"80",
          4481 => x"53",
          4482 => x"06",
          4483 => x"f8",
          4484 => x"1b",
          4485 => x"06",
          4486 => x"7b",
          4487 => x"80",
          4488 => x"2e",
          4489 => x"ff",
          4490 => x"39",
          4491 => x"e8",
          4492 => x"38",
          4493 => x"08",
          4494 => x"38",
          4495 => x"8f",
          4496 => x"c5",
          4497 => x"98",
          4498 => x"70",
          4499 => x"59",
          4500 => x"ee",
          4501 => x"ff",
          4502 => x"c4",
          4503 => x"2b",
          4504 => x"82",
          4505 => x"70",
          4506 => x"97",
          4507 => x"2c",
          4508 => x"29",
          4509 => x"05",
          4510 => x"70",
          4511 => x"51",
          4512 => x"51",
          4513 => x"81",
          4514 => x"2e",
          4515 => x"77",
          4516 => x"38",
          4517 => x"0a",
          4518 => x"0a",
          4519 => x"2c",
          4520 => x"75",
          4521 => x"38",
          4522 => x"52",
          4523 => x"85",
          4524 => x"98",
          4525 => x"06",
          4526 => x"2e",
          4527 => x"82",
          4528 => x"81",
          4529 => x"74",
          4530 => x"29",
          4531 => x"05",
          4532 => x"70",
          4533 => x"56",
          4534 => x"95",
          4535 => x"76",
          4536 => x"77",
          4537 => x"3f",
          4538 => x"08",
          4539 => x"54",
          4540 => x"d3",
          4541 => x"75",
          4542 => x"ca",
          4543 => x"55",
          4544 => x"c4",
          4545 => x"2b",
          4546 => x"82",
          4547 => x"70",
          4548 => x"98",
          4549 => x"11",
          4550 => x"82",
          4551 => x"33",
          4552 => x"51",
          4553 => x"55",
          4554 => x"09",
          4555 => x"92",
          4556 => x"ac",
          4557 => x"0c",
          4558 => x"cd",
          4559 => x"0b",
          4560 => x"34",
          4561 => x"82",
          4562 => x"75",
          4563 => x"34",
          4564 => x"34",
          4565 => x"7e",
          4566 => x"26",
          4567 => x"73",
          4568 => x"96",
          4569 => x"73",
          4570 => x"cd",
          4571 => x"73",
          4572 => x"cb",
          4573 => x"c8",
          4574 => x"75",
          4575 => x"74",
          4576 => x"98",
          4577 => x"73",
          4578 => x"38",
          4579 => x"73",
          4580 => x"34",
          4581 => x"0a",
          4582 => x"0a",
          4583 => x"2c",
          4584 => x"33",
          4585 => x"df",
          4586 => x"cc",
          4587 => x"56",
          4588 => x"cd",
          4589 => x"1a",
          4590 => x"33",
          4591 => x"cd",
          4592 => x"73",
          4593 => x"38",
          4594 => x"73",
          4595 => x"34",
          4596 => x"33",
          4597 => x"0a",
          4598 => x"0a",
          4599 => x"2c",
          4600 => x"33",
          4601 => x"56",
          4602 => x"a8",
          4603 => x"ec",
          4604 => x"1a",
          4605 => x"54",
          4606 => x"3f",
          4607 => x"0a",
          4608 => x"0a",
          4609 => x"2c",
          4610 => x"33",
          4611 => x"73",
          4612 => x"38",
          4613 => x"33",
          4614 => x"70",
          4615 => x"cd",
          4616 => x"51",
          4617 => x"77",
          4618 => x"38",
          4619 => x"08",
          4620 => x"ff",
          4621 => x"74",
          4622 => x"29",
          4623 => x"05",
          4624 => x"82",
          4625 => x"56",
          4626 => x"75",
          4627 => x"fb",
          4628 => x"7a",
          4629 => x"81",
          4630 => x"cd",
          4631 => x"52",
          4632 => x"51",
          4633 => x"81",
          4634 => x"cd",
          4635 => x"81",
          4636 => x"55",
          4637 => x"fb",
          4638 => x"cd",
          4639 => x"05",
          4640 => x"cd",
          4641 => x"15",
          4642 => x"cd",
          4643 => x"cd",
          4644 => x"88",
          4645 => x"9d",
          4646 => x"cc",
          4647 => x"2b",
          4648 => x"82",
          4649 => x"57",
          4650 => x"74",
          4651 => x"38",
          4652 => x"81",
          4653 => x"34",
          4654 => x"08",
          4655 => x"51",
          4656 => x"3f",
          4657 => x"0a",
          4658 => x"0a",
          4659 => x"2c",
          4660 => x"33",
          4661 => x"75",
          4662 => x"38",
          4663 => x"08",
          4664 => x"ff",
          4665 => x"82",
          4666 => x"70",
          4667 => x"98",
          4668 => x"c8",
          4669 => x"56",
          4670 => x"24",
          4671 => x"82",
          4672 => x"52",
          4673 => x"a1",
          4674 => x"81",
          4675 => x"81",
          4676 => x"70",
          4677 => x"cd",
          4678 => x"51",
          4679 => x"25",
          4680 => x"9b",
          4681 => x"c8",
          4682 => x"54",
          4683 => x"82",
          4684 => x"52",
          4685 => x"a0",
          4686 => x"cd",
          4687 => x"51",
          4688 => x"82",
          4689 => x"81",
          4690 => x"73",
          4691 => x"cd",
          4692 => x"73",
          4693 => x"38",
          4694 => x"52",
          4695 => x"f3",
          4696 => x"80",
          4697 => x"0b",
          4698 => x"34",
          4699 => x"cd",
          4700 => x"82",
          4701 => x"af",
          4702 => x"82",
          4703 => x"54",
          4704 => x"f9",
          4705 => x"cd",
          4706 => x"88",
          4707 => x"a5",
          4708 => x"cc",
          4709 => x"54",
          4710 => x"cc",
          4711 => x"ff",
          4712 => x"39",
          4713 => x"33",
          4714 => x"33",
          4715 => x"75",
          4716 => x"38",
          4717 => x"73",
          4718 => x"34",
          4719 => x"70",
          4720 => x"81",
          4721 => x"51",
          4722 => x"25",
          4723 => x"1a",
          4724 => x"33",
          4725 => x"cd",
          4726 => x"73",
          4727 => x"9f",
          4728 => x"81",
          4729 => x"81",
          4730 => x"70",
          4731 => x"cd",
          4732 => x"51",
          4733 => x"24",
          4734 => x"cd",
          4735 => x"a0",
          4736 => x"b1",
          4737 => x"cc",
          4738 => x"2b",
          4739 => x"82",
          4740 => x"57",
          4741 => x"74",
          4742 => x"a3",
          4743 => x"ec",
          4744 => x"51",
          4745 => x"3f",
          4746 => x"0a",
          4747 => x"0a",
          4748 => x"2c",
          4749 => x"33",
          4750 => x"75",
          4751 => x"38",
          4752 => x"82",
          4753 => x"70",
          4754 => x"82",
          4755 => x"59",
          4756 => x"77",
          4757 => x"38",
          4758 => x"08",
          4759 => x"54",
          4760 => x"cc",
          4761 => x"70",
          4762 => x"ff",
          4763 => x"82",
          4764 => x"70",
          4765 => x"82",
          4766 => x"58",
          4767 => x"75",
          4768 => x"f7",
          4769 => x"cd",
          4770 => x"52",
          4771 => x"51",
          4772 => x"80",
          4773 => x"cc",
          4774 => x"82",
          4775 => x"f7",
          4776 => x"b0",
          4777 => x"e4",
          4778 => x"80",
          4779 => x"74",
          4780 => x"d4",
          4781 => x"98",
          4782 => x"c8",
          4783 => x"98",
          4784 => x"06",
          4785 => x"74",
          4786 => x"ff",
          4787 => x"93",
          4788 => x"39",
          4789 => x"82",
          4790 => x"fc",
          4791 => x"54",
          4792 => x"a7",
          4793 => x"ff",
          4794 => x"82",
          4795 => x"82",
          4796 => x"82",
          4797 => x"81",
          4798 => x"05",
          4799 => x"79",
          4800 => x"e4",
          4801 => x"54",
          4802 => x"73",
          4803 => x"80",
          4804 => x"38",
          4805 => x"a5",
          4806 => x"39",
          4807 => x"09",
          4808 => x"38",
          4809 => x"08",
          4810 => x"2e",
          4811 => x"51",
          4812 => x"3f",
          4813 => x"08",
          4814 => x"34",
          4815 => x"08",
          4816 => x"81",
          4817 => x"52",
          4818 => x"a7",
          4819 => x"c3",
          4820 => x"29",
          4821 => x"05",
          4822 => x"54",
          4823 => x"ab",
          4824 => x"ff",
          4825 => x"82",
          4826 => x"82",
          4827 => x"82",
          4828 => x"81",
          4829 => x"05",
          4830 => x"79",
          4831 => x"e8",
          4832 => x"54",
          4833 => x"06",
          4834 => x"74",
          4835 => x"34",
          4836 => x"82",
          4837 => x"82",
          4838 => x"52",
          4839 => x"e2",
          4840 => x"39",
          4841 => x"33",
          4842 => x"06",
          4843 => x"33",
          4844 => x"74",
          4845 => x"87",
          4846 => x"ec",
          4847 => x"14",
          4848 => x"cd",
          4849 => x"1a",
          4850 => x"54",
          4851 => x"3f",
          4852 => x"82",
          4853 => x"54",
          4854 => x"f4",
          4855 => x"cd",
          4856 => x"88",
          4857 => x"cd",
          4858 => x"cc",
          4859 => x"54",
          4860 => x"cc",
          4861 => x"39",
          4862 => x"83",
          4863 => x"82",
          4864 => x"84",
          4865 => x"b6",
          4866 => x"80",
          4867 => x"83",
          4868 => x"ff",
          4869 => x"82",
          4870 => x"54",
          4871 => x"74",
          4872 => x"76",
          4873 => x"82",
          4874 => x"54",
          4875 => x"34",
          4876 => x"34",
          4877 => x"08",
          4878 => x"15",
          4879 => x"15",
          4880 => x"90",
          4881 => x"8c",
          4882 => x"fe",
          4883 => x"70",
          4884 => x"06",
          4885 => x"58",
          4886 => x"74",
          4887 => x"73",
          4888 => x"82",
          4889 => x"70",
          4890 => x"b6",
          4891 => x"f8",
          4892 => x"55",
          4893 => x"34",
          4894 => x"34",
          4895 => x"04",
          4896 => x"73",
          4897 => x"84",
          4898 => x"38",
          4899 => x"2a",
          4900 => x"83",
          4901 => x"51",
          4902 => x"82",
          4903 => x"83",
          4904 => x"f9",
          4905 => x"a6",
          4906 => x"84",
          4907 => x"22",
          4908 => x"b6",
          4909 => x"83",
          4910 => x"74",
          4911 => x"11",
          4912 => x"12",
          4913 => x"2b",
          4914 => x"05",
          4915 => x"71",
          4916 => x"06",
          4917 => x"2a",
          4918 => x"59",
          4919 => x"57",
          4920 => x"71",
          4921 => x"81",
          4922 => x"b6",
          4923 => x"75",
          4924 => x"54",
          4925 => x"34",
          4926 => x"34",
          4927 => x"08",
          4928 => x"33",
          4929 => x"71",
          4930 => x"70",
          4931 => x"ff",
          4932 => x"52",
          4933 => x"05",
          4934 => x"ff",
          4935 => x"2a",
          4936 => x"71",
          4937 => x"72",
          4938 => x"53",
          4939 => x"34",
          4940 => x"08",
          4941 => x"76",
          4942 => x"17",
          4943 => x"0d",
          4944 => x"0d",
          4945 => x"08",
          4946 => x"9e",
          4947 => x"83",
          4948 => x"86",
          4949 => x"12",
          4950 => x"2b",
          4951 => x"07",
          4952 => x"52",
          4953 => x"05",
          4954 => x"85",
          4955 => x"88",
          4956 => x"88",
          4957 => x"56",
          4958 => x"13",
          4959 => x"13",
          4960 => x"90",
          4961 => x"84",
          4962 => x"12",
          4963 => x"2b",
          4964 => x"07",
          4965 => x"52",
          4966 => x"12",
          4967 => x"33",
          4968 => x"07",
          4969 => x"54",
          4970 => x"70",
          4971 => x"73",
          4972 => x"82",
          4973 => x"13",
          4974 => x"12",
          4975 => x"2b",
          4976 => x"ff",
          4977 => x"88",
          4978 => x"53",
          4979 => x"73",
          4980 => x"14",
          4981 => x"0d",
          4982 => x"0d",
          4983 => x"22",
          4984 => x"08",
          4985 => x"71",
          4986 => x"81",
          4987 => x"88",
          4988 => x"88",
          4989 => x"33",
          4990 => x"71",
          4991 => x"90",
          4992 => x"5f",
          4993 => x"5a",
          4994 => x"54",
          4995 => x"80",
          4996 => x"51",
          4997 => x"82",
          4998 => x"70",
          4999 => x"81",
          5000 => x"8b",
          5001 => x"2b",
          5002 => x"70",
          5003 => x"33",
          5004 => x"07",
          5005 => x"8f",
          5006 => x"51",
          5007 => x"53",
          5008 => x"72",
          5009 => x"2a",
          5010 => x"82",
          5011 => x"83",
          5012 => x"b6",
          5013 => x"16",
          5014 => x"12",
          5015 => x"2b",
          5016 => x"07",
          5017 => x"55",
          5018 => x"33",
          5019 => x"71",
          5020 => x"70",
          5021 => x"06",
          5022 => x"57",
          5023 => x"52",
          5024 => x"71",
          5025 => x"88",
          5026 => x"fb",
          5027 => x"b6",
          5028 => x"84",
          5029 => x"22",
          5030 => x"72",
          5031 => x"33",
          5032 => x"71",
          5033 => x"83",
          5034 => x"5b",
          5035 => x"52",
          5036 => x"33",
          5037 => x"71",
          5038 => x"02",
          5039 => x"05",
          5040 => x"70",
          5041 => x"51",
          5042 => x"71",
          5043 => x"81",
          5044 => x"b6",
          5045 => x"15",
          5046 => x"12",
          5047 => x"2b",
          5048 => x"07",
          5049 => x"52",
          5050 => x"12",
          5051 => x"33",
          5052 => x"07",
          5053 => x"54",
          5054 => x"70",
          5055 => x"72",
          5056 => x"82",
          5057 => x"14",
          5058 => x"83",
          5059 => x"88",
          5060 => x"b6",
          5061 => x"54",
          5062 => x"04",
          5063 => x"7b",
          5064 => x"08",
          5065 => x"70",
          5066 => x"06",
          5067 => x"53",
          5068 => x"82",
          5069 => x"76",
          5070 => x"11",
          5071 => x"83",
          5072 => x"8b",
          5073 => x"2b",
          5074 => x"70",
          5075 => x"33",
          5076 => x"71",
          5077 => x"53",
          5078 => x"53",
          5079 => x"59",
          5080 => x"25",
          5081 => x"80",
          5082 => x"51",
          5083 => x"81",
          5084 => x"14",
          5085 => x"33",
          5086 => x"71",
          5087 => x"76",
          5088 => x"2a",
          5089 => x"58",
          5090 => x"14",
          5091 => x"ff",
          5092 => x"87",
          5093 => x"b6",
          5094 => x"19",
          5095 => x"85",
          5096 => x"88",
          5097 => x"88",
          5098 => x"5b",
          5099 => x"84",
          5100 => x"85",
          5101 => x"b6",
          5102 => x"53",
          5103 => x"14",
          5104 => x"87",
          5105 => x"b6",
          5106 => x"76",
          5107 => x"75",
          5108 => x"82",
          5109 => x"18",
          5110 => x"12",
          5111 => x"2b",
          5112 => x"80",
          5113 => x"88",
          5114 => x"55",
          5115 => x"74",
          5116 => x"15",
          5117 => x"0d",
          5118 => x"0d",
          5119 => x"b6",
          5120 => x"38",
          5121 => x"71",
          5122 => x"38",
          5123 => x"8c",
          5124 => x"0d",
          5125 => x"0d",
          5126 => x"58",
          5127 => x"82",
          5128 => x"83",
          5129 => x"82",
          5130 => x"84",
          5131 => x"12",
          5132 => x"2b",
          5133 => x"59",
          5134 => x"81",
          5135 => x"75",
          5136 => x"cb",
          5137 => x"29",
          5138 => x"81",
          5139 => x"88",
          5140 => x"81",
          5141 => x"79",
          5142 => x"ff",
          5143 => x"7f",
          5144 => x"51",
          5145 => x"77",
          5146 => x"38",
          5147 => x"85",
          5148 => x"5a",
          5149 => x"33",
          5150 => x"71",
          5151 => x"57",
          5152 => x"38",
          5153 => x"ff",
          5154 => x"7a",
          5155 => x"80",
          5156 => x"82",
          5157 => x"11",
          5158 => x"12",
          5159 => x"2b",
          5160 => x"ff",
          5161 => x"52",
          5162 => x"55",
          5163 => x"83",
          5164 => x"80",
          5165 => x"26",
          5166 => x"74",
          5167 => x"2e",
          5168 => x"77",
          5169 => x"81",
          5170 => x"75",
          5171 => x"3f",
          5172 => x"82",
          5173 => x"79",
          5174 => x"f7",
          5175 => x"b6",
          5176 => x"1c",
          5177 => x"87",
          5178 => x"8b",
          5179 => x"2b",
          5180 => x"5e",
          5181 => x"7a",
          5182 => x"ff",
          5183 => x"88",
          5184 => x"56",
          5185 => x"15",
          5186 => x"ff",
          5187 => x"85",
          5188 => x"b6",
          5189 => x"83",
          5190 => x"72",
          5191 => x"33",
          5192 => x"71",
          5193 => x"70",
          5194 => x"5b",
          5195 => x"56",
          5196 => x"19",
          5197 => x"19",
          5198 => x"90",
          5199 => x"84",
          5200 => x"12",
          5201 => x"2b",
          5202 => x"07",
          5203 => x"55",
          5204 => x"78",
          5205 => x"76",
          5206 => x"82",
          5207 => x"70",
          5208 => x"84",
          5209 => x"12",
          5210 => x"2b",
          5211 => x"2a",
          5212 => x"52",
          5213 => x"84",
          5214 => x"85",
          5215 => x"b6",
          5216 => x"84",
          5217 => x"82",
          5218 => x"8d",
          5219 => x"fe",
          5220 => x"52",
          5221 => x"08",
          5222 => x"dc",
          5223 => x"71",
          5224 => x"38",
          5225 => x"ed",
          5226 => x"98",
          5227 => x"82",
          5228 => x"84",
          5229 => x"ee",
          5230 => x"66",
          5231 => x"70",
          5232 => x"b6",
          5233 => x"2e",
          5234 => x"84",
          5235 => x"3f",
          5236 => x"7e",
          5237 => x"3f",
          5238 => x"08",
          5239 => x"39",
          5240 => x"7b",
          5241 => x"3f",
          5242 => x"ba",
          5243 => x"f5",
          5244 => x"b6",
          5245 => x"ff",
          5246 => x"b6",
          5247 => x"71",
          5248 => x"70",
          5249 => x"06",
          5250 => x"73",
          5251 => x"81",
          5252 => x"88",
          5253 => x"75",
          5254 => x"ff",
          5255 => x"88",
          5256 => x"73",
          5257 => x"70",
          5258 => x"33",
          5259 => x"07",
          5260 => x"53",
          5261 => x"48",
          5262 => x"54",
          5263 => x"56",
          5264 => x"80",
          5265 => x"76",
          5266 => x"06",
          5267 => x"83",
          5268 => x"42",
          5269 => x"33",
          5270 => x"71",
          5271 => x"70",
          5272 => x"70",
          5273 => x"33",
          5274 => x"71",
          5275 => x"53",
          5276 => x"56",
          5277 => x"25",
          5278 => x"75",
          5279 => x"ff",
          5280 => x"54",
          5281 => x"81",
          5282 => x"18",
          5283 => x"2e",
          5284 => x"8f",
          5285 => x"f6",
          5286 => x"83",
          5287 => x"58",
          5288 => x"7f",
          5289 => x"74",
          5290 => x"78",
          5291 => x"3f",
          5292 => x"7f",
          5293 => x"75",
          5294 => x"38",
          5295 => x"11",
          5296 => x"33",
          5297 => x"07",
          5298 => x"f4",
          5299 => x"52",
          5300 => x"b7",
          5301 => x"98",
          5302 => x"ff",
          5303 => x"7c",
          5304 => x"2b",
          5305 => x"08",
          5306 => x"53",
          5307 => x"93",
          5308 => x"b6",
          5309 => x"84",
          5310 => x"ff",
          5311 => x"5c",
          5312 => x"60",
          5313 => x"74",
          5314 => x"38",
          5315 => x"c9",
          5316 => x"90",
          5317 => x"11",
          5318 => x"33",
          5319 => x"07",
          5320 => x"f4",
          5321 => x"52",
          5322 => x"df",
          5323 => x"98",
          5324 => x"ff",
          5325 => x"7c",
          5326 => x"2b",
          5327 => x"08",
          5328 => x"53",
          5329 => x"92",
          5330 => x"b6",
          5331 => x"84",
          5332 => x"05",
          5333 => x"73",
          5334 => x"06",
          5335 => x"7b",
          5336 => x"f9",
          5337 => x"b6",
          5338 => x"82",
          5339 => x"80",
          5340 => x"7d",
          5341 => x"82",
          5342 => x"51",
          5343 => x"3f",
          5344 => x"98",
          5345 => x"7a",
          5346 => x"38",
          5347 => x"52",
          5348 => x"8f",
          5349 => x"83",
          5350 => x"90",
          5351 => x"05",
          5352 => x"3f",
          5353 => x"82",
          5354 => x"94",
          5355 => x"fc",
          5356 => x"77",
          5357 => x"54",
          5358 => x"82",
          5359 => x"55",
          5360 => x"08",
          5361 => x"38",
          5362 => x"52",
          5363 => x"08",
          5364 => x"95",
          5365 => x"b6",
          5366 => x"3d",
          5367 => x"3d",
          5368 => x"05",
          5369 => x"52",
          5370 => x"87",
          5371 => x"94",
          5372 => x"71",
          5373 => x"0c",
          5374 => x"04",
          5375 => x"02",
          5376 => x"02",
          5377 => x"05",
          5378 => x"83",
          5379 => x"26",
          5380 => x"72",
          5381 => x"c0",
          5382 => x"53",
          5383 => x"74",
          5384 => x"38",
          5385 => x"73",
          5386 => x"c0",
          5387 => x"51",
          5388 => x"85",
          5389 => x"98",
          5390 => x"52",
          5391 => x"82",
          5392 => x"70",
          5393 => x"38",
          5394 => x"8c",
          5395 => x"ec",
          5396 => x"fc",
          5397 => x"52",
          5398 => x"87",
          5399 => x"08",
          5400 => x"2e",
          5401 => x"82",
          5402 => x"34",
          5403 => x"13",
          5404 => x"82",
          5405 => x"86",
          5406 => x"f3",
          5407 => x"62",
          5408 => x"05",
          5409 => x"57",
          5410 => x"83",
          5411 => x"fe",
          5412 => x"b6",
          5413 => x"06",
          5414 => x"71",
          5415 => x"71",
          5416 => x"2b",
          5417 => x"80",
          5418 => x"92",
          5419 => x"c0",
          5420 => x"41",
          5421 => x"5a",
          5422 => x"87",
          5423 => x"0c",
          5424 => x"84",
          5425 => x"08",
          5426 => x"70",
          5427 => x"53",
          5428 => x"2e",
          5429 => x"08",
          5430 => x"70",
          5431 => x"34",
          5432 => x"80",
          5433 => x"53",
          5434 => x"2e",
          5435 => x"53",
          5436 => x"26",
          5437 => x"80",
          5438 => x"87",
          5439 => x"08",
          5440 => x"38",
          5441 => x"8c",
          5442 => x"80",
          5443 => x"78",
          5444 => x"99",
          5445 => x"0c",
          5446 => x"8c",
          5447 => x"08",
          5448 => x"51",
          5449 => x"38",
          5450 => x"8d",
          5451 => x"17",
          5452 => x"81",
          5453 => x"53",
          5454 => x"2e",
          5455 => x"fc",
          5456 => x"52",
          5457 => x"7d",
          5458 => x"ed",
          5459 => x"80",
          5460 => x"71",
          5461 => x"38",
          5462 => x"53",
          5463 => x"98",
          5464 => x"0d",
          5465 => x"0d",
          5466 => x"02",
          5467 => x"05",
          5468 => x"58",
          5469 => x"80",
          5470 => x"fc",
          5471 => x"b6",
          5472 => x"06",
          5473 => x"71",
          5474 => x"81",
          5475 => x"38",
          5476 => x"2b",
          5477 => x"80",
          5478 => x"92",
          5479 => x"c0",
          5480 => x"40",
          5481 => x"5a",
          5482 => x"c0",
          5483 => x"76",
          5484 => x"76",
          5485 => x"75",
          5486 => x"2a",
          5487 => x"51",
          5488 => x"80",
          5489 => x"7a",
          5490 => x"5c",
          5491 => x"81",
          5492 => x"81",
          5493 => x"06",
          5494 => x"80",
          5495 => x"87",
          5496 => x"08",
          5497 => x"38",
          5498 => x"8c",
          5499 => x"80",
          5500 => x"77",
          5501 => x"99",
          5502 => x"0c",
          5503 => x"8c",
          5504 => x"08",
          5505 => x"51",
          5506 => x"38",
          5507 => x"8d",
          5508 => x"70",
          5509 => x"84",
          5510 => x"5b",
          5511 => x"2e",
          5512 => x"fc",
          5513 => x"52",
          5514 => x"7d",
          5515 => x"f8",
          5516 => x"80",
          5517 => x"71",
          5518 => x"38",
          5519 => x"53",
          5520 => x"98",
          5521 => x"0d",
          5522 => x"0d",
          5523 => x"05",
          5524 => x"02",
          5525 => x"05",
          5526 => x"54",
          5527 => x"fe",
          5528 => x"98",
          5529 => x"53",
          5530 => x"80",
          5531 => x"0b",
          5532 => x"8c",
          5533 => x"71",
          5534 => x"dc",
          5535 => x"24",
          5536 => x"84",
          5537 => x"92",
          5538 => x"54",
          5539 => x"8d",
          5540 => x"39",
          5541 => x"80",
          5542 => x"cb",
          5543 => x"70",
          5544 => x"81",
          5545 => x"52",
          5546 => x"8a",
          5547 => x"98",
          5548 => x"71",
          5549 => x"c0",
          5550 => x"52",
          5551 => x"81",
          5552 => x"c0",
          5553 => x"53",
          5554 => x"82",
          5555 => x"71",
          5556 => x"39",
          5557 => x"39",
          5558 => x"77",
          5559 => x"81",
          5560 => x"72",
          5561 => x"84",
          5562 => x"73",
          5563 => x"0c",
          5564 => x"04",
          5565 => x"74",
          5566 => x"71",
          5567 => x"2b",
          5568 => x"98",
          5569 => x"84",
          5570 => x"fd",
          5571 => x"83",
          5572 => x"12",
          5573 => x"2b",
          5574 => x"07",
          5575 => x"70",
          5576 => x"2b",
          5577 => x"07",
          5578 => x"0c",
          5579 => x"56",
          5580 => x"3d",
          5581 => x"3d",
          5582 => x"84",
          5583 => x"22",
          5584 => x"72",
          5585 => x"54",
          5586 => x"2a",
          5587 => x"34",
          5588 => x"04",
          5589 => x"73",
          5590 => x"70",
          5591 => x"05",
          5592 => x"88",
          5593 => x"72",
          5594 => x"54",
          5595 => x"2a",
          5596 => x"70",
          5597 => x"34",
          5598 => x"51",
          5599 => x"83",
          5600 => x"fe",
          5601 => x"75",
          5602 => x"51",
          5603 => x"92",
          5604 => x"81",
          5605 => x"73",
          5606 => x"55",
          5607 => x"51",
          5608 => x"3d",
          5609 => x"3d",
          5610 => x"76",
          5611 => x"72",
          5612 => x"05",
          5613 => x"11",
          5614 => x"38",
          5615 => x"04",
          5616 => x"78",
          5617 => x"56",
          5618 => x"81",
          5619 => x"74",
          5620 => x"56",
          5621 => x"31",
          5622 => x"52",
          5623 => x"80",
          5624 => x"71",
          5625 => x"38",
          5626 => x"98",
          5627 => x"0d",
          5628 => x"0d",
          5629 => x"51",
          5630 => x"73",
          5631 => x"81",
          5632 => x"33",
          5633 => x"38",
          5634 => x"b6",
          5635 => x"3d",
          5636 => x"0b",
          5637 => x"0c",
          5638 => x"82",
          5639 => x"04",
          5640 => x"7b",
          5641 => x"83",
          5642 => x"5a",
          5643 => x"80",
          5644 => x"54",
          5645 => x"53",
          5646 => x"53",
          5647 => x"52",
          5648 => x"3f",
          5649 => x"08",
          5650 => x"81",
          5651 => x"82",
          5652 => x"83",
          5653 => x"16",
          5654 => x"18",
          5655 => x"18",
          5656 => x"58",
          5657 => x"9f",
          5658 => x"33",
          5659 => x"2e",
          5660 => x"93",
          5661 => x"76",
          5662 => x"52",
          5663 => x"51",
          5664 => x"83",
          5665 => x"79",
          5666 => x"0c",
          5667 => x"04",
          5668 => x"78",
          5669 => x"80",
          5670 => x"17",
          5671 => x"38",
          5672 => x"fc",
          5673 => x"98",
          5674 => x"b6",
          5675 => x"38",
          5676 => x"53",
          5677 => x"81",
          5678 => x"f7",
          5679 => x"b6",
          5680 => x"2e",
          5681 => x"55",
          5682 => x"b0",
          5683 => x"82",
          5684 => x"88",
          5685 => x"f8",
          5686 => x"70",
          5687 => x"c0",
          5688 => x"98",
          5689 => x"b6",
          5690 => x"91",
          5691 => x"55",
          5692 => x"09",
          5693 => x"f0",
          5694 => x"33",
          5695 => x"2e",
          5696 => x"80",
          5697 => x"80",
          5698 => x"98",
          5699 => x"17",
          5700 => x"fd",
          5701 => x"d4",
          5702 => x"b2",
          5703 => x"96",
          5704 => x"85",
          5705 => x"75",
          5706 => x"3f",
          5707 => x"e4",
          5708 => x"98",
          5709 => x"9c",
          5710 => x"08",
          5711 => x"17",
          5712 => x"3f",
          5713 => x"52",
          5714 => x"51",
          5715 => x"a0",
          5716 => x"05",
          5717 => x"0c",
          5718 => x"75",
          5719 => x"33",
          5720 => x"3f",
          5721 => x"34",
          5722 => x"52",
          5723 => x"51",
          5724 => x"82",
          5725 => x"80",
          5726 => x"81",
          5727 => x"b6",
          5728 => x"3d",
          5729 => x"3d",
          5730 => x"1a",
          5731 => x"fe",
          5732 => x"54",
          5733 => x"73",
          5734 => x"8a",
          5735 => x"71",
          5736 => x"08",
          5737 => x"75",
          5738 => x"0c",
          5739 => x"04",
          5740 => x"7a",
          5741 => x"56",
          5742 => x"77",
          5743 => x"38",
          5744 => x"08",
          5745 => x"38",
          5746 => x"54",
          5747 => x"2e",
          5748 => x"72",
          5749 => x"38",
          5750 => x"8d",
          5751 => x"39",
          5752 => x"81",
          5753 => x"b6",
          5754 => x"2a",
          5755 => x"2a",
          5756 => x"05",
          5757 => x"55",
          5758 => x"82",
          5759 => x"81",
          5760 => x"83",
          5761 => x"b4",
          5762 => x"17",
          5763 => x"a4",
          5764 => x"55",
          5765 => x"57",
          5766 => x"3f",
          5767 => x"08",
          5768 => x"74",
          5769 => x"14",
          5770 => x"70",
          5771 => x"07",
          5772 => x"71",
          5773 => x"52",
          5774 => x"72",
          5775 => x"75",
          5776 => x"58",
          5777 => x"76",
          5778 => x"15",
          5779 => x"73",
          5780 => x"3f",
          5781 => x"08",
          5782 => x"76",
          5783 => x"06",
          5784 => x"05",
          5785 => x"3f",
          5786 => x"08",
          5787 => x"06",
          5788 => x"76",
          5789 => x"15",
          5790 => x"73",
          5791 => x"3f",
          5792 => x"08",
          5793 => x"82",
          5794 => x"06",
          5795 => x"05",
          5796 => x"3f",
          5797 => x"08",
          5798 => x"58",
          5799 => x"58",
          5800 => x"98",
          5801 => x"0d",
          5802 => x"0d",
          5803 => x"5a",
          5804 => x"59",
          5805 => x"82",
          5806 => x"98",
          5807 => x"82",
          5808 => x"33",
          5809 => x"2e",
          5810 => x"72",
          5811 => x"38",
          5812 => x"8d",
          5813 => x"39",
          5814 => x"81",
          5815 => x"f7",
          5816 => x"2a",
          5817 => x"2a",
          5818 => x"05",
          5819 => x"55",
          5820 => x"82",
          5821 => x"59",
          5822 => x"08",
          5823 => x"74",
          5824 => x"16",
          5825 => x"16",
          5826 => x"59",
          5827 => x"53",
          5828 => x"8f",
          5829 => x"2b",
          5830 => x"74",
          5831 => x"71",
          5832 => x"72",
          5833 => x"0b",
          5834 => x"74",
          5835 => x"17",
          5836 => x"75",
          5837 => x"3f",
          5838 => x"08",
          5839 => x"98",
          5840 => x"38",
          5841 => x"06",
          5842 => x"78",
          5843 => x"54",
          5844 => x"77",
          5845 => x"33",
          5846 => x"71",
          5847 => x"51",
          5848 => x"34",
          5849 => x"76",
          5850 => x"17",
          5851 => x"75",
          5852 => x"3f",
          5853 => x"08",
          5854 => x"98",
          5855 => x"38",
          5856 => x"ff",
          5857 => x"10",
          5858 => x"76",
          5859 => x"51",
          5860 => x"be",
          5861 => x"2a",
          5862 => x"05",
          5863 => x"f9",
          5864 => x"b6",
          5865 => x"82",
          5866 => x"ab",
          5867 => x"0a",
          5868 => x"2b",
          5869 => x"70",
          5870 => x"70",
          5871 => x"54",
          5872 => x"82",
          5873 => x"8f",
          5874 => x"07",
          5875 => x"f7",
          5876 => x"0b",
          5877 => x"78",
          5878 => x"0c",
          5879 => x"04",
          5880 => x"7a",
          5881 => x"08",
          5882 => x"59",
          5883 => x"a4",
          5884 => x"17",
          5885 => x"38",
          5886 => x"aa",
          5887 => x"73",
          5888 => x"fd",
          5889 => x"b6",
          5890 => x"82",
          5891 => x"80",
          5892 => x"39",
          5893 => x"eb",
          5894 => x"80",
          5895 => x"b6",
          5896 => x"80",
          5897 => x"52",
          5898 => x"84",
          5899 => x"98",
          5900 => x"b6",
          5901 => x"2e",
          5902 => x"82",
          5903 => x"81",
          5904 => x"82",
          5905 => x"ff",
          5906 => x"80",
          5907 => x"75",
          5908 => x"3f",
          5909 => x"08",
          5910 => x"16",
          5911 => x"90",
          5912 => x"55",
          5913 => x"27",
          5914 => x"15",
          5915 => x"84",
          5916 => x"07",
          5917 => x"17",
          5918 => x"76",
          5919 => x"a6",
          5920 => x"73",
          5921 => x"0c",
          5922 => x"04",
          5923 => x"7c",
          5924 => x"59",
          5925 => x"95",
          5926 => x"08",
          5927 => x"2e",
          5928 => x"17",
          5929 => x"b2",
          5930 => x"ae",
          5931 => x"7a",
          5932 => x"3f",
          5933 => x"82",
          5934 => x"27",
          5935 => x"82",
          5936 => x"55",
          5937 => x"08",
          5938 => x"d2",
          5939 => x"08",
          5940 => x"08",
          5941 => x"38",
          5942 => x"17",
          5943 => x"54",
          5944 => x"82",
          5945 => x"7a",
          5946 => x"06",
          5947 => x"81",
          5948 => x"17",
          5949 => x"83",
          5950 => x"75",
          5951 => x"f9",
          5952 => x"59",
          5953 => x"08",
          5954 => x"81",
          5955 => x"82",
          5956 => x"59",
          5957 => x"08",
          5958 => x"70",
          5959 => x"25",
          5960 => x"82",
          5961 => x"54",
          5962 => x"55",
          5963 => x"38",
          5964 => x"08",
          5965 => x"38",
          5966 => x"54",
          5967 => x"90",
          5968 => x"18",
          5969 => x"38",
          5970 => x"39",
          5971 => x"38",
          5972 => x"16",
          5973 => x"08",
          5974 => x"38",
          5975 => x"78",
          5976 => x"38",
          5977 => x"51",
          5978 => x"82",
          5979 => x"80",
          5980 => x"80",
          5981 => x"98",
          5982 => x"09",
          5983 => x"38",
          5984 => x"08",
          5985 => x"98",
          5986 => x"30",
          5987 => x"80",
          5988 => x"07",
          5989 => x"55",
          5990 => x"38",
          5991 => x"09",
          5992 => x"ae",
          5993 => x"80",
          5994 => x"53",
          5995 => x"51",
          5996 => x"82",
          5997 => x"82",
          5998 => x"30",
          5999 => x"98",
          6000 => x"25",
          6001 => x"79",
          6002 => x"38",
          6003 => x"8f",
          6004 => x"79",
          6005 => x"f9",
          6006 => x"b6",
          6007 => x"74",
          6008 => x"8c",
          6009 => x"17",
          6010 => x"90",
          6011 => x"54",
          6012 => x"86",
          6013 => x"90",
          6014 => x"17",
          6015 => x"54",
          6016 => x"34",
          6017 => x"56",
          6018 => x"90",
          6019 => x"80",
          6020 => x"82",
          6021 => x"55",
          6022 => x"56",
          6023 => x"82",
          6024 => x"8c",
          6025 => x"f8",
          6026 => x"70",
          6027 => x"f0",
          6028 => x"98",
          6029 => x"56",
          6030 => x"08",
          6031 => x"7b",
          6032 => x"f6",
          6033 => x"b6",
          6034 => x"b6",
          6035 => x"17",
          6036 => x"80",
          6037 => x"b4",
          6038 => x"57",
          6039 => x"77",
          6040 => x"81",
          6041 => x"15",
          6042 => x"78",
          6043 => x"81",
          6044 => x"53",
          6045 => x"15",
          6046 => x"e9",
          6047 => x"98",
          6048 => x"df",
          6049 => x"22",
          6050 => x"30",
          6051 => x"70",
          6052 => x"51",
          6053 => x"82",
          6054 => x"8a",
          6055 => x"f8",
          6056 => x"7c",
          6057 => x"56",
          6058 => x"80",
          6059 => x"f1",
          6060 => x"06",
          6061 => x"e9",
          6062 => x"18",
          6063 => x"08",
          6064 => x"38",
          6065 => x"82",
          6066 => x"38",
          6067 => x"54",
          6068 => x"74",
          6069 => x"82",
          6070 => x"22",
          6071 => x"79",
          6072 => x"38",
          6073 => x"98",
          6074 => x"cd",
          6075 => x"22",
          6076 => x"54",
          6077 => x"26",
          6078 => x"52",
          6079 => x"b0",
          6080 => x"98",
          6081 => x"b6",
          6082 => x"2e",
          6083 => x"0b",
          6084 => x"08",
          6085 => x"98",
          6086 => x"b6",
          6087 => x"85",
          6088 => x"bd",
          6089 => x"31",
          6090 => x"73",
          6091 => x"f4",
          6092 => x"b6",
          6093 => x"18",
          6094 => x"18",
          6095 => x"08",
          6096 => x"72",
          6097 => x"38",
          6098 => x"58",
          6099 => x"89",
          6100 => x"18",
          6101 => x"ff",
          6102 => x"05",
          6103 => x"80",
          6104 => x"b6",
          6105 => x"3d",
          6106 => x"3d",
          6107 => x"08",
          6108 => x"a0",
          6109 => x"54",
          6110 => x"77",
          6111 => x"80",
          6112 => x"0c",
          6113 => x"53",
          6114 => x"80",
          6115 => x"38",
          6116 => x"06",
          6117 => x"b5",
          6118 => x"98",
          6119 => x"14",
          6120 => x"92",
          6121 => x"2a",
          6122 => x"56",
          6123 => x"26",
          6124 => x"80",
          6125 => x"16",
          6126 => x"77",
          6127 => x"53",
          6128 => x"38",
          6129 => x"51",
          6130 => x"82",
          6131 => x"53",
          6132 => x"0b",
          6133 => x"08",
          6134 => x"38",
          6135 => x"b6",
          6136 => x"2e",
          6137 => x"98",
          6138 => x"b6",
          6139 => x"80",
          6140 => x"8a",
          6141 => x"15",
          6142 => x"80",
          6143 => x"14",
          6144 => x"51",
          6145 => x"82",
          6146 => x"53",
          6147 => x"b6",
          6148 => x"2e",
          6149 => x"82",
          6150 => x"98",
          6151 => x"ba",
          6152 => x"82",
          6153 => x"ff",
          6154 => x"82",
          6155 => x"52",
          6156 => x"f3",
          6157 => x"98",
          6158 => x"72",
          6159 => x"72",
          6160 => x"f2",
          6161 => x"b6",
          6162 => x"15",
          6163 => x"15",
          6164 => x"b4",
          6165 => x"0c",
          6166 => x"82",
          6167 => x"8a",
          6168 => x"f7",
          6169 => x"7d",
          6170 => x"5b",
          6171 => x"76",
          6172 => x"3f",
          6173 => x"08",
          6174 => x"98",
          6175 => x"38",
          6176 => x"08",
          6177 => x"08",
          6178 => x"f0",
          6179 => x"b6",
          6180 => x"82",
          6181 => x"80",
          6182 => x"b6",
          6183 => x"18",
          6184 => x"51",
          6185 => x"81",
          6186 => x"81",
          6187 => x"81",
          6188 => x"98",
          6189 => x"83",
          6190 => x"77",
          6191 => x"72",
          6192 => x"38",
          6193 => x"75",
          6194 => x"81",
          6195 => x"a5",
          6196 => x"98",
          6197 => x"52",
          6198 => x"8e",
          6199 => x"98",
          6200 => x"b6",
          6201 => x"2e",
          6202 => x"73",
          6203 => x"81",
          6204 => x"87",
          6205 => x"b6",
          6206 => x"3d",
          6207 => x"3d",
          6208 => x"11",
          6209 => x"ec",
          6210 => x"98",
          6211 => x"ff",
          6212 => x"33",
          6213 => x"71",
          6214 => x"81",
          6215 => x"94",
          6216 => x"d0",
          6217 => x"98",
          6218 => x"73",
          6219 => x"82",
          6220 => x"85",
          6221 => x"fc",
          6222 => x"79",
          6223 => x"ff",
          6224 => x"12",
          6225 => x"eb",
          6226 => x"70",
          6227 => x"72",
          6228 => x"81",
          6229 => x"73",
          6230 => x"94",
          6231 => x"d6",
          6232 => x"0d",
          6233 => x"0d",
          6234 => x"55",
          6235 => x"5a",
          6236 => x"08",
          6237 => x"8a",
          6238 => x"08",
          6239 => x"ee",
          6240 => x"b6",
          6241 => x"82",
          6242 => x"80",
          6243 => x"15",
          6244 => x"55",
          6245 => x"38",
          6246 => x"e6",
          6247 => x"33",
          6248 => x"70",
          6249 => x"58",
          6250 => x"86",
          6251 => x"b6",
          6252 => x"73",
          6253 => x"83",
          6254 => x"73",
          6255 => x"38",
          6256 => x"06",
          6257 => x"80",
          6258 => x"75",
          6259 => x"38",
          6260 => x"08",
          6261 => x"54",
          6262 => x"2e",
          6263 => x"83",
          6264 => x"73",
          6265 => x"38",
          6266 => x"51",
          6267 => x"82",
          6268 => x"58",
          6269 => x"08",
          6270 => x"15",
          6271 => x"38",
          6272 => x"0b",
          6273 => x"77",
          6274 => x"0c",
          6275 => x"04",
          6276 => x"77",
          6277 => x"54",
          6278 => x"51",
          6279 => x"82",
          6280 => x"55",
          6281 => x"08",
          6282 => x"14",
          6283 => x"51",
          6284 => x"82",
          6285 => x"55",
          6286 => x"08",
          6287 => x"53",
          6288 => x"08",
          6289 => x"08",
          6290 => x"3f",
          6291 => x"14",
          6292 => x"08",
          6293 => x"3f",
          6294 => x"17",
          6295 => x"b6",
          6296 => x"3d",
          6297 => x"3d",
          6298 => x"08",
          6299 => x"54",
          6300 => x"53",
          6301 => x"82",
          6302 => x"8d",
          6303 => x"08",
          6304 => x"34",
          6305 => x"15",
          6306 => x"0d",
          6307 => x"0d",
          6308 => x"57",
          6309 => x"17",
          6310 => x"08",
          6311 => x"82",
          6312 => x"89",
          6313 => x"55",
          6314 => x"14",
          6315 => x"16",
          6316 => x"71",
          6317 => x"38",
          6318 => x"09",
          6319 => x"38",
          6320 => x"73",
          6321 => x"81",
          6322 => x"ae",
          6323 => x"05",
          6324 => x"15",
          6325 => x"70",
          6326 => x"34",
          6327 => x"8a",
          6328 => x"38",
          6329 => x"05",
          6330 => x"81",
          6331 => x"17",
          6332 => x"12",
          6333 => x"34",
          6334 => x"9c",
          6335 => x"e8",
          6336 => x"b6",
          6337 => x"0c",
          6338 => x"e7",
          6339 => x"b6",
          6340 => x"17",
          6341 => x"51",
          6342 => x"82",
          6343 => x"84",
          6344 => x"3d",
          6345 => x"3d",
          6346 => x"08",
          6347 => x"61",
          6348 => x"55",
          6349 => x"2e",
          6350 => x"55",
          6351 => x"2e",
          6352 => x"80",
          6353 => x"94",
          6354 => x"1c",
          6355 => x"81",
          6356 => x"61",
          6357 => x"56",
          6358 => x"2e",
          6359 => x"83",
          6360 => x"73",
          6361 => x"70",
          6362 => x"25",
          6363 => x"51",
          6364 => x"38",
          6365 => x"0c",
          6366 => x"51",
          6367 => x"26",
          6368 => x"80",
          6369 => x"34",
          6370 => x"51",
          6371 => x"82",
          6372 => x"55",
          6373 => x"91",
          6374 => x"1d",
          6375 => x"8b",
          6376 => x"79",
          6377 => x"3f",
          6378 => x"57",
          6379 => x"55",
          6380 => x"2e",
          6381 => x"80",
          6382 => x"18",
          6383 => x"1a",
          6384 => x"70",
          6385 => x"2a",
          6386 => x"07",
          6387 => x"5a",
          6388 => x"8c",
          6389 => x"54",
          6390 => x"81",
          6391 => x"39",
          6392 => x"70",
          6393 => x"2a",
          6394 => x"75",
          6395 => x"8c",
          6396 => x"2e",
          6397 => x"a0",
          6398 => x"38",
          6399 => x"0c",
          6400 => x"76",
          6401 => x"38",
          6402 => x"b8",
          6403 => x"70",
          6404 => x"5a",
          6405 => x"76",
          6406 => x"38",
          6407 => x"70",
          6408 => x"dc",
          6409 => x"72",
          6410 => x"80",
          6411 => x"51",
          6412 => x"73",
          6413 => x"38",
          6414 => x"18",
          6415 => x"1a",
          6416 => x"55",
          6417 => x"2e",
          6418 => x"83",
          6419 => x"73",
          6420 => x"70",
          6421 => x"25",
          6422 => x"51",
          6423 => x"38",
          6424 => x"75",
          6425 => x"81",
          6426 => x"81",
          6427 => x"27",
          6428 => x"73",
          6429 => x"38",
          6430 => x"70",
          6431 => x"32",
          6432 => x"80",
          6433 => x"2a",
          6434 => x"56",
          6435 => x"81",
          6436 => x"57",
          6437 => x"f5",
          6438 => x"2b",
          6439 => x"25",
          6440 => x"80",
          6441 => x"af",
          6442 => x"57",
          6443 => x"e6",
          6444 => x"b6",
          6445 => x"2e",
          6446 => x"18",
          6447 => x"1a",
          6448 => x"56",
          6449 => x"3f",
          6450 => x"08",
          6451 => x"e8",
          6452 => x"54",
          6453 => x"80",
          6454 => x"17",
          6455 => x"34",
          6456 => x"11",
          6457 => x"74",
          6458 => x"75",
          6459 => x"80",
          6460 => x"3f",
          6461 => x"08",
          6462 => x"9f",
          6463 => x"99",
          6464 => x"e0",
          6465 => x"ff",
          6466 => x"79",
          6467 => x"74",
          6468 => x"57",
          6469 => x"77",
          6470 => x"76",
          6471 => x"38",
          6472 => x"73",
          6473 => x"09",
          6474 => x"38",
          6475 => x"84",
          6476 => x"27",
          6477 => x"39",
          6478 => x"f2",
          6479 => x"80",
          6480 => x"54",
          6481 => x"34",
          6482 => x"58",
          6483 => x"f2",
          6484 => x"b6",
          6485 => x"82",
          6486 => x"80",
          6487 => x"1b",
          6488 => x"51",
          6489 => x"82",
          6490 => x"56",
          6491 => x"08",
          6492 => x"9c",
          6493 => x"33",
          6494 => x"80",
          6495 => x"38",
          6496 => x"bf",
          6497 => x"86",
          6498 => x"15",
          6499 => x"2a",
          6500 => x"51",
          6501 => x"92",
          6502 => x"79",
          6503 => x"e4",
          6504 => x"b6",
          6505 => x"2e",
          6506 => x"52",
          6507 => x"ba",
          6508 => x"39",
          6509 => x"33",
          6510 => x"80",
          6511 => x"74",
          6512 => x"81",
          6513 => x"38",
          6514 => x"70",
          6515 => x"82",
          6516 => x"54",
          6517 => x"96",
          6518 => x"06",
          6519 => x"2e",
          6520 => x"ff",
          6521 => x"1c",
          6522 => x"80",
          6523 => x"81",
          6524 => x"ba",
          6525 => x"b6",
          6526 => x"2a",
          6527 => x"51",
          6528 => x"38",
          6529 => x"70",
          6530 => x"81",
          6531 => x"55",
          6532 => x"e1",
          6533 => x"08",
          6534 => x"1d",
          6535 => x"7c",
          6536 => x"3f",
          6537 => x"08",
          6538 => x"fa",
          6539 => x"82",
          6540 => x"8f",
          6541 => x"f6",
          6542 => x"5b",
          6543 => x"70",
          6544 => x"59",
          6545 => x"73",
          6546 => x"c6",
          6547 => x"81",
          6548 => x"70",
          6549 => x"52",
          6550 => x"8d",
          6551 => x"38",
          6552 => x"09",
          6553 => x"a5",
          6554 => x"d0",
          6555 => x"ff",
          6556 => x"53",
          6557 => x"91",
          6558 => x"73",
          6559 => x"d0",
          6560 => x"71",
          6561 => x"f7",
          6562 => x"82",
          6563 => x"55",
          6564 => x"55",
          6565 => x"81",
          6566 => x"74",
          6567 => x"56",
          6568 => x"12",
          6569 => x"70",
          6570 => x"38",
          6571 => x"81",
          6572 => x"51",
          6573 => x"51",
          6574 => x"89",
          6575 => x"70",
          6576 => x"53",
          6577 => x"70",
          6578 => x"51",
          6579 => x"09",
          6580 => x"38",
          6581 => x"38",
          6582 => x"77",
          6583 => x"70",
          6584 => x"2a",
          6585 => x"07",
          6586 => x"51",
          6587 => x"8f",
          6588 => x"84",
          6589 => x"83",
          6590 => x"94",
          6591 => x"74",
          6592 => x"38",
          6593 => x"0c",
          6594 => x"86",
          6595 => x"e4",
          6596 => x"82",
          6597 => x"8c",
          6598 => x"fa",
          6599 => x"56",
          6600 => x"17",
          6601 => x"b0",
          6602 => x"52",
          6603 => x"e0",
          6604 => x"82",
          6605 => x"81",
          6606 => x"b2",
          6607 => x"b4",
          6608 => x"98",
          6609 => x"ff",
          6610 => x"55",
          6611 => x"d5",
          6612 => x"06",
          6613 => x"80",
          6614 => x"33",
          6615 => x"81",
          6616 => x"81",
          6617 => x"81",
          6618 => x"eb",
          6619 => x"70",
          6620 => x"07",
          6621 => x"73",
          6622 => x"81",
          6623 => x"81",
          6624 => x"83",
          6625 => x"90",
          6626 => x"16",
          6627 => x"3f",
          6628 => x"08",
          6629 => x"98",
          6630 => x"9d",
          6631 => x"82",
          6632 => x"81",
          6633 => x"e0",
          6634 => x"b6",
          6635 => x"82",
          6636 => x"80",
          6637 => x"82",
          6638 => x"b6",
          6639 => x"3d",
          6640 => x"3d",
          6641 => x"84",
          6642 => x"05",
          6643 => x"80",
          6644 => x"51",
          6645 => x"82",
          6646 => x"58",
          6647 => x"0b",
          6648 => x"08",
          6649 => x"38",
          6650 => x"08",
          6651 => x"cd",
          6652 => x"08",
          6653 => x"56",
          6654 => x"86",
          6655 => x"75",
          6656 => x"fe",
          6657 => x"54",
          6658 => x"2e",
          6659 => x"14",
          6660 => x"ca",
          6661 => x"98",
          6662 => x"06",
          6663 => x"54",
          6664 => x"38",
          6665 => x"86",
          6666 => x"82",
          6667 => x"06",
          6668 => x"56",
          6669 => x"38",
          6670 => x"80",
          6671 => x"81",
          6672 => x"52",
          6673 => x"51",
          6674 => x"82",
          6675 => x"81",
          6676 => x"81",
          6677 => x"83",
          6678 => x"87",
          6679 => x"2e",
          6680 => x"82",
          6681 => x"06",
          6682 => x"56",
          6683 => x"38",
          6684 => x"74",
          6685 => x"a3",
          6686 => x"98",
          6687 => x"06",
          6688 => x"2e",
          6689 => x"80",
          6690 => x"3d",
          6691 => x"83",
          6692 => x"15",
          6693 => x"53",
          6694 => x"8d",
          6695 => x"15",
          6696 => x"3f",
          6697 => x"08",
          6698 => x"70",
          6699 => x"0c",
          6700 => x"16",
          6701 => x"80",
          6702 => x"80",
          6703 => x"54",
          6704 => x"84",
          6705 => x"5b",
          6706 => x"80",
          6707 => x"7a",
          6708 => x"fc",
          6709 => x"b6",
          6710 => x"ff",
          6711 => x"77",
          6712 => x"81",
          6713 => x"76",
          6714 => x"81",
          6715 => x"2e",
          6716 => x"8d",
          6717 => x"26",
          6718 => x"bf",
          6719 => x"f4",
          6720 => x"98",
          6721 => x"ff",
          6722 => x"84",
          6723 => x"81",
          6724 => x"38",
          6725 => x"51",
          6726 => x"82",
          6727 => x"83",
          6728 => x"58",
          6729 => x"80",
          6730 => x"db",
          6731 => x"b6",
          6732 => x"77",
          6733 => x"80",
          6734 => x"82",
          6735 => x"c4",
          6736 => x"11",
          6737 => x"06",
          6738 => x"8d",
          6739 => x"26",
          6740 => x"74",
          6741 => x"78",
          6742 => x"c1",
          6743 => x"59",
          6744 => x"15",
          6745 => x"2e",
          6746 => x"13",
          6747 => x"72",
          6748 => x"38",
          6749 => x"eb",
          6750 => x"14",
          6751 => x"3f",
          6752 => x"08",
          6753 => x"98",
          6754 => x"23",
          6755 => x"57",
          6756 => x"83",
          6757 => x"c7",
          6758 => x"d8",
          6759 => x"98",
          6760 => x"ff",
          6761 => x"8d",
          6762 => x"14",
          6763 => x"3f",
          6764 => x"08",
          6765 => x"14",
          6766 => x"3f",
          6767 => x"08",
          6768 => x"06",
          6769 => x"72",
          6770 => x"97",
          6771 => x"22",
          6772 => x"84",
          6773 => x"5a",
          6774 => x"83",
          6775 => x"14",
          6776 => x"79",
          6777 => x"f3",
          6778 => x"b6",
          6779 => x"82",
          6780 => x"80",
          6781 => x"38",
          6782 => x"08",
          6783 => x"ff",
          6784 => x"38",
          6785 => x"83",
          6786 => x"83",
          6787 => x"74",
          6788 => x"85",
          6789 => x"89",
          6790 => x"76",
          6791 => x"c3",
          6792 => x"70",
          6793 => x"7b",
          6794 => x"73",
          6795 => x"17",
          6796 => x"ac",
          6797 => x"55",
          6798 => x"09",
          6799 => x"38",
          6800 => x"51",
          6801 => x"82",
          6802 => x"83",
          6803 => x"53",
          6804 => x"82",
          6805 => x"82",
          6806 => x"e0",
          6807 => x"ab",
          6808 => x"98",
          6809 => x"0c",
          6810 => x"53",
          6811 => x"56",
          6812 => x"81",
          6813 => x"13",
          6814 => x"74",
          6815 => x"82",
          6816 => x"74",
          6817 => x"81",
          6818 => x"06",
          6819 => x"83",
          6820 => x"2a",
          6821 => x"72",
          6822 => x"26",
          6823 => x"ff",
          6824 => x"0c",
          6825 => x"15",
          6826 => x"0b",
          6827 => x"76",
          6828 => x"81",
          6829 => x"38",
          6830 => x"51",
          6831 => x"82",
          6832 => x"83",
          6833 => x"53",
          6834 => x"09",
          6835 => x"f9",
          6836 => x"52",
          6837 => x"b8",
          6838 => x"98",
          6839 => x"38",
          6840 => x"08",
          6841 => x"84",
          6842 => x"d8",
          6843 => x"b6",
          6844 => x"ff",
          6845 => x"72",
          6846 => x"2e",
          6847 => x"80",
          6848 => x"14",
          6849 => x"3f",
          6850 => x"08",
          6851 => x"a4",
          6852 => x"81",
          6853 => x"84",
          6854 => x"d7",
          6855 => x"b6",
          6856 => x"8a",
          6857 => x"2e",
          6858 => x"9d",
          6859 => x"14",
          6860 => x"3f",
          6861 => x"08",
          6862 => x"84",
          6863 => x"d7",
          6864 => x"b6",
          6865 => x"15",
          6866 => x"34",
          6867 => x"22",
          6868 => x"72",
          6869 => x"23",
          6870 => x"23",
          6871 => x"15",
          6872 => x"75",
          6873 => x"0c",
          6874 => x"04",
          6875 => x"77",
          6876 => x"73",
          6877 => x"38",
          6878 => x"72",
          6879 => x"38",
          6880 => x"71",
          6881 => x"38",
          6882 => x"84",
          6883 => x"52",
          6884 => x"09",
          6885 => x"38",
          6886 => x"51",
          6887 => x"82",
          6888 => x"81",
          6889 => x"88",
          6890 => x"08",
          6891 => x"39",
          6892 => x"73",
          6893 => x"74",
          6894 => x"0c",
          6895 => x"04",
          6896 => x"02",
          6897 => x"7a",
          6898 => x"fc",
          6899 => x"f4",
          6900 => x"54",
          6901 => x"b6",
          6902 => x"bc",
          6903 => x"98",
          6904 => x"82",
          6905 => x"70",
          6906 => x"73",
          6907 => x"38",
          6908 => x"78",
          6909 => x"2e",
          6910 => x"74",
          6911 => x"0c",
          6912 => x"80",
          6913 => x"80",
          6914 => x"70",
          6915 => x"51",
          6916 => x"82",
          6917 => x"54",
          6918 => x"98",
          6919 => x"0d",
          6920 => x"0d",
          6921 => x"05",
          6922 => x"33",
          6923 => x"54",
          6924 => x"84",
          6925 => x"bf",
          6926 => x"98",
          6927 => x"53",
          6928 => x"05",
          6929 => x"fa",
          6930 => x"98",
          6931 => x"b6",
          6932 => x"a4",
          6933 => x"68",
          6934 => x"70",
          6935 => x"c6",
          6936 => x"98",
          6937 => x"b6",
          6938 => x"38",
          6939 => x"05",
          6940 => x"2b",
          6941 => x"80",
          6942 => x"86",
          6943 => x"06",
          6944 => x"2e",
          6945 => x"74",
          6946 => x"38",
          6947 => x"09",
          6948 => x"38",
          6949 => x"f8",
          6950 => x"98",
          6951 => x"39",
          6952 => x"33",
          6953 => x"73",
          6954 => x"77",
          6955 => x"81",
          6956 => x"73",
          6957 => x"38",
          6958 => x"bc",
          6959 => x"07",
          6960 => x"b4",
          6961 => x"2a",
          6962 => x"51",
          6963 => x"2e",
          6964 => x"62",
          6965 => x"e8",
          6966 => x"b6",
          6967 => x"82",
          6968 => x"52",
          6969 => x"51",
          6970 => x"62",
          6971 => x"8b",
          6972 => x"53",
          6973 => x"51",
          6974 => x"80",
          6975 => x"05",
          6976 => x"3f",
          6977 => x"0b",
          6978 => x"75",
          6979 => x"f1",
          6980 => x"11",
          6981 => x"80",
          6982 => x"97",
          6983 => x"51",
          6984 => x"82",
          6985 => x"55",
          6986 => x"08",
          6987 => x"b7",
          6988 => x"c4",
          6989 => x"05",
          6990 => x"2a",
          6991 => x"51",
          6992 => x"80",
          6993 => x"84",
          6994 => x"39",
          6995 => x"70",
          6996 => x"54",
          6997 => x"a9",
          6998 => x"06",
          6999 => x"2e",
          7000 => x"55",
          7001 => x"73",
          7002 => x"d6",
          7003 => x"b6",
          7004 => x"ff",
          7005 => x"0c",
          7006 => x"b6",
          7007 => x"f8",
          7008 => x"2a",
          7009 => x"51",
          7010 => x"2e",
          7011 => x"80",
          7012 => x"7a",
          7013 => x"a0",
          7014 => x"a4",
          7015 => x"53",
          7016 => x"e6",
          7017 => x"b6",
          7018 => x"b6",
          7019 => x"1b",
          7020 => x"05",
          7021 => x"d3",
          7022 => x"98",
          7023 => x"98",
          7024 => x"0c",
          7025 => x"56",
          7026 => x"84",
          7027 => x"90",
          7028 => x"0b",
          7029 => x"80",
          7030 => x"0c",
          7031 => x"1a",
          7032 => x"2a",
          7033 => x"51",
          7034 => x"2e",
          7035 => x"82",
          7036 => x"80",
          7037 => x"38",
          7038 => x"08",
          7039 => x"8a",
          7040 => x"89",
          7041 => x"59",
          7042 => x"76",
          7043 => x"d7",
          7044 => x"b6",
          7045 => x"82",
          7046 => x"81",
          7047 => x"82",
          7048 => x"98",
          7049 => x"09",
          7050 => x"38",
          7051 => x"78",
          7052 => x"30",
          7053 => x"80",
          7054 => x"77",
          7055 => x"38",
          7056 => x"06",
          7057 => x"c3",
          7058 => x"1a",
          7059 => x"38",
          7060 => x"06",
          7061 => x"2e",
          7062 => x"52",
          7063 => x"a6",
          7064 => x"98",
          7065 => x"82",
          7066 => x"75",
          7067 => x"b6",
          7068 => x"9c",
          7069 => x"39",
          7070 => x"74",
          7071 => x"b6",
          7072 => x"3d",
          7073 => x"3d",
          7074 => x"65",
          7075 => x"5d",
          7076 => x"0c",
          7077 => x"05",
          7078 => x"f9",
          7079 => x"b6",
          7080 => x"82",
          7081 => x"8a",
          7082 => x"33",
          7083 => x"2e",
          7084 => x"56",
          7085 => x"90",
          7086 => x"06",
          7087 => x"74",
          7088 => x"b6",
          7089 => x"82",
          7090 => x"34",
          7091 => x"aa",
          7092 => x"91",
          7093 => x"56",
          7094 => x"8c",
          7095 => x"1a",
          7096 => x"74",
          7097 => x"38",
          7098 => x"80",
          7099 => x"38",
          7100 => x"70",
          7101 => x"56",
          7102 => x"b2",
          7103 => x"11",
          7104 => x"77",
          7105 => x"5b",
          7106 => x"38",
          7107 => x"88",
          7108 => x"8f",
          7109 => x"08",
          7110 => x"d5",
          7111 => x"b6",
          7112 => x"81",
          7113 => x"9f",
          7114 => x"2e",
          7115 => x"74",
          7116 => x"98",
          7117 => x"7e",
          7118 => x"3f",
          7119 => x"08",
          7120 => x"83",
          7121 => x"98",
          7122 => x"89",
          7123 => x"77",
          7124 => x"d6",
          7125 => x"7f",
          7126 => x"58",
          7127 => x"75",
          7128 => x"75",
          7129 => x"77",
          7130 => x"7c",
          7131 => x"33",
          7132 => x"3f",
          7133 => x"08",
          7134 => x"7e",
          7135 => x"56",
          7136 => x"2e",
          7137 => x"16",
          7138 => x"55",
          7139 => x"94",
          7140 => x"53",
          7141 => x"b0",
          7142 => x"31",
          7143 => x"05",
          7144 => x"3f",
          7145 => x"56",
          7146 => x"9c",
          7147 => x"19",
          7148 => x"06",
          7149 => x"31",
          7150 => x"76",
          7151 => x"7b",
          7152 => x"08",
          7153 => x"d1",
          7154 => x"b6",
          7155 => x"81",
          7156 => x"94",
          7157 => x"ff",
          7158 => x"05",
          7159 => x"cf",
          7160 => x"76",
          7161 => x"17",
          7162 => x"1e",
          7163 => x"18",
          7164 => x"5e",
          7165 => x"39",
          7166 => x"82",
          7167 => x"90",
          7168 => x"f2",
          7169 => x"63",
          7170 => x"40",
          7171 => x"7e",
          7172 => x"fc",
          7173 => x"51",
          7174 => x"82",
          7175 => x"55",
          7176 => x"08",
          7177 => x"18",
          7178 => x"80",
          7179 => x"74",
          7180 => x"39",
          7181 => x"70",
          7182 => x"81",
          7183 => x"56",
          7184 => x"80",
          7185 => x"38",
          7186 => x"0b",
          7187 => x"82",
          7188 => x"39",
          7189 => x"19",
          7190 => x"83",
          7191 => x"18",
          7192 => x"56",
          7193 => x"27",
          7194 => x"09",
          7195 => x"2e",
          7196 => x"94",
          7197 => x"83",
          7198 => x"56",
          7199 => x"38",
          7200 => x"22",
          7201 => x"89",
          7202 => x"55",
          7203 => x"75",
          7204 => x"18",
          7205 => x"9c",
          7206 => x"85",
          7207 => x"08",
          7208 => x"d7",
          7209 => x"b6",
          7210 => x"82",
          7211 => x"80",
          7212 => x"38",
          7213 => x"ff",
          7214 => x"ff",
          7215 => x"38",
          7216 => x"0c",
          7217 => x"85",
          7218 => x"19",
          7219 => x"b0",
          7220 => x"19",
          7221 => x"81",
          7222 => x"74",
          7223 => x"3f",
          7224 => x"08",
          7225 => x"98",
          7226 => x"7e",
          7227 => x"3f",
          7228 => x"08",
          7229 => x"d2",
          7230 => x"98",
          7231 => x"89",
          7232 => x"78",
          7233 => x"d5",
          7234 => x"7f",
          7235 => x"58",
          7236 => x"75",
          7237 => x"75",
          7238 => x"78",
          7239 => x"7c",
          7240 => x"33",
          7241 => x"3f",
          7242 => x"08",
          7243 => x"7e",
          7244 => x"78",
          7245 => x"74",
          7246 => x"38",
          7247 => x"b0",
          7248 => x"31",
          7249 => x"05",
          7250 => x"51",
          7251 => x"7e",
          7252 => x"83",
          7253 => x"89",
          7254 => x"db",
          7255 => x"08",
          7256 => x"26",
          7257 => x"51",
          7258 => x"82",
          7259 => x"fd",
          7260 => x"77",
          7261 => x"55",
          7262 => x"0c",
          7263 => x"83",
          7264 => x"80",
          7265 => x"55",
          7266 => x"83",
          7267 => x"9c",
          7268 => x"7e",
          7269 => x"3f",
          7270 => x"08",
          7271 => x"75",
          7272 => x"94",
          7273 => x"ff",
          7274 => x"05",
          7275 => x"3f",
          7276 => x"0b",
          7277 => x"7b",
          7278 => x"08",
          7279 => x"76",
          7280 => x"08",
          7281 => x"1c",
          7282 => x"08",
          7283 => x"5c",
          7284 => x"83",
          7285 => x"74",
          7286 => x"fd",
          7287 => x"18",
          7288 => x"07",
          7289 => x"19",
          7290 => x"75",
          7291 => x"0c",
          7292 => x"04",
          7293 => x"7a",
          7294 => x"05",
          7295 => x"56",
          7296 => x"82",
          7297 => x"57",
          7298 => x"08",
          7299 => x"90",
          7300 => x"86",
          7301 => x"06",
          7302 => x"73",
          7303 => x"e9",
          7304 => x"08",
          7305 => x"cc",
          7306 => x"b6",
          7307 => x"82",
          7308 => x"80",
          7309 => x"16",
          7310 => x"33",
          7311 => x"55",
          7312 => x"34",
          7313 => x"53",
          7314 => x"08",
          7315 => x"3f",
          7316 => x"52",
          7317 => x"c9",
          7318 => x"88",
          7319 => x"96",
          7320 => x"f0",
          7321 => x"92",
          7322 => x"ca",
          7323 => x"81",
          7324 => x"34",
          7325 => x"df",
          7326 => x"98",
          7327 => x"33",
          7328 => x"55",
          7329 => x"17",
          7330 => x"b6",
          7331 => x"3d",
          7332 => x"3d",
          7333 => x"52",
          7334 => x"3f",
          7335 => x"08",
          7336 => x"98",
          7337 => x"86",
          7338 => x"52",
          7339 => x"bc",
          7340 => x"98",
          7341 => x"b6",
          7342 => x"38",
          7343 => x"08",
          7344 => x"82",
          7345 => x"86",
          7346 => x"ff",
          7347 => x"3d",
          7348 => x"3f",
          7349 => x"0b",
          7350 => x"08",
          7351 => x"82",
          7352 => x"82",
          7353 => x"80",
          7354 => x"b6",
          7355 => x"3d",
          7356 => x"3d",
          7357 => x"93",
          7358 => x"52",
          7359 => x"e9",
          7360 => x"b6",
          7361 => x"82",
          7362 => x"80",
          7363 => x"58",
          7364 => x"3d",
          7365 => x"e0",
          7366 => x"b6",
          7367 => x"82",
          7368 => x"bc",
          7369 => x"c7",
          7370 => x"98",
          7371 => x"73",
          7372 => x"38",
          7373 => x"12",
          7374 => x"39",
          7375 => x"33",
          7376 => x"70",
          7377 => x"55",
          7378 => x"2e",
          7379 => x"7f",
          7380 => x"54",
          7381 => x"82",
          7382 => x"94",
          7383 => x"39",
          7384 => x"08",
          7385 => x"81",
          7386 => x"85",
          7387 => x"b6",
          7388 => x"3d",
          7389 => x"3d",
          7390 => x"5b",
          7391 => x"34",
          7392 => x"3d",
          7393 => x"52",
          7394 => x"e8",
          7395 => x"b6",
          7396 => x"82",
          7397 => x"82",
          7398 => x"43",
          7399 => x"11",
          7400 => x"58",
          7401 => x"80",
          7402 => x"38",
          7403 => x"3d",
          7404 => x"d5",
          7405 => x"b6",
          7406 => x"82",
          7407 => x"82",
          7408 => x"52",
          7409 => x"c8",
          7410 => x"98",
          7411 => x"b6",
          7412 => x"c1",
          7413 => x"7b",
          7414 => x"3f",
          7415 => x"08",
          7416 => x"74",
          7417 => x"3f",
          7418 => x"08",
          7419 => x"98",
          7420 => x"38",
          7421 => x"51",
          7422 => x"82",
          7423 => x"57",
          7424 => x"08",
          7425 => x"52",
          7426 => x"f2",
          7427 => x"b6",
          7428 => x"a6",
          7429 => x"74",
          7430 => x"3f",
          7431 => x"08",
          7432 => x"98",
          7433 => x"cc",
          7434 => x"2e",
          7435 => x"86",
          7436 => x"81",
          7437 => x"81",
          7438 => x"3d",
          7439 => x"52",
          7440 => x"c9",
          7441 => x"3d",
          7442 => x"11",
          7443 => x"5a",
          7444 => x"2e",
          7445 => x"b9",
          7446 => x"16",
          7447 => x"33",
          7448 => x"73",
          7449 => x"16",
          7450 => x"26",
          7451 => x"75",
          7452 => x"38",
          7453 => x"05",
          7454 => x"6f",
          7455 => x"ff",
          7456 => x"55",
          7457 => x"74",
          7458 => x"38",
          7459 => x"11",
          7460 => x"74",
          7461 => x"39",
          7462 => x"09",
          7463 => x"38",
          7464 => x"11",
          7465 => x"74",
          7466 => x"82",
          7467 => x"70",
          7468 => x"af",
          7469 => x"08",
          7470 => x"5c",
          7471 => x"73",
          7472 => x"38",
          7473 => x"1a",
          7474 => x"55",
          7475 => x"38",
          7476 => x"73",
          7477 => x"38",
          7478 => x"76",
          7479 => x"74",
          7480 => x"33",
          7481 => x"05",
          7482 => x"15",
          7483 => x"ba",
          7484 => x"05",
          7485 => x"ff",
          7486 => x"06",
          7487 => x"57",
          7488 => x"18",
          7489 => x"54",
          7490 => x"70",
          7491 => x"34",
          7492 => x"ee",
          7493 => x"34",
          7494 => x"98",
          7495 => x"0d",
          7496 => x"0d",
          7497 => x"3d",
          7498 => x"71",
          7499 => x"ec",
          7500 => x"b6",
          7501 => x"82",
          7502 => x"82",
          7503 => x"15",
          7504 => x"82",
          7505 => x"15",
          7506 => x"76",
          7507 => x"90",
          7508 => x"81",
          7509 => x"06",
          7510 => x"72",
          7511 => x"56",
          7512 => x"54",
          7513 => x"17",
          7514 => x"78",
          7515 => x"38",
          7516 => x"22",
          7517 => x"59",
          7518 => x"78",
          7519 => x"76",
          7520 => x"51",
          7521 => x"3f",
          7522 => x"08",
          7523 => x"54",
          7524 => x"53",
          7525 => x"3f",
          7526 => x"08",
          7527 => x"38",
          7528 => x"75",
          7529 => x"18",
          7530 => x"31",
          7531 => x"57",
          7532 => x"b1",
          7533 => x"08",
          7534 => x"38",
          7535 => x"51",
          7536 => x"82",
          7537 => x"54",
          7538 => x"08",
          7539 => x"9a",
          7540 => x"98",
          7541 => x"81",
          7542 => x"b6",
          7543 => x"16",
          7544 => x"16",
          7545 => x"2e",
          7546 => x"76",
          7547 => x"dc",
          7548 => x"31",
          7549 => x"18",
          7550 => x"90",
          7551 => x"81",
          7552 => x"06",
          7553 => x"56",
          7554 => x"9a",
          7555 => x"74",
          7556 => x"3f",
          7557 => x"08",
          7558 => x"98",
          7559 => x"82",
          7560 => x"56",
          7561 => x"52",
          7562 => x"84",
          7563 => x"98",
          7564 => x"ff",
          7565 => x"81",
          7566 => x"38",
          7567 => x"98",
          7568 => x"a6",
          7569 => x"16",
          7570 => x"39",
          7571 => x"16",
          7572 => x"75",
          7573 => x"53",
          7574 => x"aa",
          7575 => x"79",
          7576 => x"3f",
          7577 => x"08",
          7578 => x"0b",
          7579 => x"82",
          7580 => x"39",
          7581 => x"16",
          7582 => x"bb",
          7583 => x"2a",
          7584 => x"08",
          7585 => x"15",
          7586 => x"15",
          7587 => x"90",
          7588 => x"16",
          7589 => x"33",
          7590 => x"53",
          7591 => x"34",
          7592 => x"06",
          7593 => x"2e",
          7594 => x"9c",
          7595 => x"85",
          7596 => x"16",
          7597 => x"72",
          7598 => x"0c",
          7599 => x"04",
          7600 => x"79",
          7601 => x"75",
          7602 => x"8a",
          7603 => x"89",
          7604 => x"52",
          7605 => x"05",
          7606 => x"3f",
          7607 => x"08",
          7608 => x"98",
          7609 => x"38",
          7610 => x"7a",
          7611 => x"d8",
          7612 => x"b6",
          7613 => x"82",
          7614 => x"80",
          7615 => x"16",
          7616 => x"2b",
          7617 => x"74",
          7618 => x"86",
          7619 => x"84",
          7620 => x"06",
          7621 => x"73",
          7622 => x"38",
          7623 => x"52",
          7624 => x"da",
          7625 => x"98",
          7626 => x"0c",
          7627 => x"14",
          7628 => x"23",
          7629 => x"51",
          7630 => x"82",
          7631 => x"55",
          7632 => x"09",
          7633 => x"38",
          7634 => x"39",
          7635 => x"84",
          7636 => x"0c",
          7637 => x"82",
          7638 => x"89",
          7639 => x"fc",
          7640 => x"87",
          7641 => x"53",
          7642 => x"e7",
          7643 => x"b6",
          7644 => x"38",
          7645 => x"08",
          7646 => x"3d",
          7647 => x"3d",
          7648 => x"89",
          7649 => x"54",
          7650 => x"54",
          7651 => x"82",
          7652 => x"53",
          7653 => x"08",
          7654 => x"74",
          7655 => x"b6",
          7656 => x"73",
          7657 => x"3f",
          7658 => x"08",
          7659 => x"39",
          7660 => x"08",
          7661 => x"d3",
          7662 => x"b6",
          7663 => x"82",
          7664 => x"84",
          7665 => x"06",
          7666 => x"53",
          7667 => x"b6",
          7668 => x"38",
          7669 => x"51",
          7670 => x"72",
          7671 => x"cf",
          7672 => x"b6",
          7673 => x"32",
          7674 => x"72",
          7675 => x"70",
          7676 => x"08",
          7677 => x"54",
          7678 => x"b6",
          7679 => x"3d",
          7680 => x"3d",
          7681 => x"80",
          7682 => x"70",
          7683 => x"52",
          7684 => x"3f",
          7685 => x"08",
          7686 => x"98",
          7687 => x"64",
          7688 => x"d6",
          7689 => x"b6",
          7690 => x"82",
          7691 => x"a0",
          7692 => x"cb",
          7693 => x"98",
          7694 => x"73",
          7695 => x"38",
          7696 => x"39",
          7697 => x"88",
          7698 => x"75",
          7699 => x"3f",
          7700 => x"98",
          7701 => x"0d",
          7702 => x"0d",
          7703 => x"5c",
          7704 => x"3d",
          7705 => x"93",
          7706 => x"d6",
          7707 => x"98",
          7708 => x"b6",
          7709 => x"80",
          7710 => x"0c",
          7711 => x"11",
          7712 => x"90",
          7713 => x"56",
          7714 => x"74",
          7715 => x"75",
          7716 => x"e4",
          7717 => x"81",
          7718 => x"5b",
          7719 => x"82",
          7720 => x"75",
          7721 => x"73",
          7722 => x"81",
          7723 => x"82",
          7724 => x"76",
          7725 => x"f0",
          7726 => x"f4",
          7727 => x"98",
          7728 => x"d1",
          7729 => x"98",
          7730 => x"ce",
          7731 => x"98",
          7732 => x"82",
          7733 => x"07",
          7734 => x"05",
          7735 => x"53",
          7736 => x"98",
          7737 => x"26",
          7738 => x"f9",
          7739 => x"08",
          7740 => x"08",
          7741 => x"98",
          7742 => x"81",
          7743 => x"58",
          7744 => x"3f",
          7745 => x"08",
          7746 => x"98",
          7747 => x"38",
          7748 => x"77",
          7749 => x"5d",
          7750 => x"74",
          7751 => x"81",
          7752 => x"b4",
          7753 => x"bb",
          7754 => x"b6",
          7755 => x"ff",
          7756 => x"30",
          7757 => x"1b",
          7758 => x"5b",
          7759 => x"39",
          7760 => x"ff",
          7761 => x"82",
          7762 => x"f0",
          7763 => x"30",
          7764 => x"1b",
          7765 => x"5b",
          7766 => x"83",
          7767 => x"58",
          7768 => x"92",
          7769 => x"0c",
          7770 => x"12",
          7771 => x"33",
          7772 => x"54",
          7773 => x"34",
          7774 => x"98",
          7775 => x"0d",
          7776 => x"0d",
          7777 => x"fc",
          7778 => x"52",
          7779 => x"3f",
          7780 => x"08",
          7781 => x"98",
          7782 => x"38",
          7783 => x"56",
          7784 => x"38",
          7785 => x"70",
          7786 => x"81",
          7787 => x"55",
          7788 => x"80",
          7789 => x"38",
          7790 => x"54",
          7791 => x"08",
          7792 => x"38",
          7793 => x"82",
          7794 => x"53",
          7795 => x"52",
          7796 => x"8c",
          7797 => x"98",
          7798 => x"19",
          7799 => x"c9",
          7800 => x"08",
          7801 => x"ff",
          7802 => x"82",
          7803 => x"ff",
          7804 => x"06",
          7805 => x"56",
          7806 => x"08",
          7807 => x"81",
          7808 => x"82",
          7809 => x"75",
          7810 => x"54",
          7811 => x"08",
          7812 => x"27",
          7813 => x"17",
          7814 => x"b6",
          7815 => x"76",
          7816 => x"3f",
          7817 => x"08",
          7818 => x"08",
          7819 => x"90",
          7820 => x"c0",
          7821 => x"90",
          7822 => x"80",
          7823 => x"75",
          7824 => x"75",
          7825 => x"b6",
          7826 => x"3d",
          7827 => x"3d",
          7828 => x"a0",
          7829 => x"05",
          7830 => x"51",
          7831 => x"82",
          7832 => x"55",
          7833 => x"08",
          7834 => x"78",
          7835 => x"08",
          7836 => x"70",
          7837 => x"ae",
          7838 => x"98",
          7839 => x"b6",
          7840 => x"db",
          7841 => x"fb",
          7842 => x"85",
          7843 => x"06",
          7844 => x"86",
          7845 => x"c7",
          7846 => x"2b",
          7847 => x"24",
          7848 => x"02",
          7849 => x"33",
          7850 => x"58",
          7851 => x"76",
          7852 => x"6b",
          7853 => x"cc",
          7854 => x"b6",
          7855 => x"84",
          7856 => x"06",
          7857 => x"73",
          7858 => x"d4",
          7859 => x"82",
          7860 => x"94",
          7861 => x"81",
          7862 => x"5a",
          7863 => x"08",
          7864 => x"8a",
          7865 => x"54",
          7866 => x"82",
          7867 => x"55",
          7868 => x"08",
          7869 => x"82",
          7870 => x"52",
          7871 => x"e5",
          7872 => x"98",
          7873 => x"b6",
          7874 => x"38",
          7875 => x"cf",
          7876 => x"98",
          7877 => x"88",
          7878 => x"98",
          7879 => x"38",
          7880 => x"c2",
          7881 => x"98",
          7882 => x"98",
          7883 => x"82",
          7884 => x"07",
          7885 => x"55",
          7886 => x"2e",
          7887 => x"80",
          7888 => x"80",
          7889 => x"77",
          7890 => x"3f",
          7891 => x"08",
          7892 => x"38",
          7893 => x"ba",
          7894 => x"b6",
          7895 => x"74",
          7896 => x"0c",
          7897 => x"04",
          7898 => x"82",
          7899 => x"c0",
          7900 => x"3d",
          7901 => x"3f",
          7902 => x"08",
          7903 => x"98",
          7904 => x"38",
          7905 => x"52",
          7906 => x"52",
          7907 => x"3f",
          7908 => x"08",
          7909 => x"98",
          7910 => x"88",
          7911 => x"39",
          7912 => x"08",
          7913 => x"81",
          7914 => x"38",
          7915 => x"05",
          7916 => x"2a",
          7917 => x"55",
          7918 => x"81",
          7919 => x"5a",
          7920 => x"3d",
          7921 => x"c1",
          7922 => x"b6",
          7923 => x"55",
          7924 => x"98",
          7925 => x"87",
          7926 => x"98",
          7927 => x"09",
          7928 => x"38",
          7929 => x"b6",
          7930 => x"2e",
          7931 => x"86",
          7932 => x"81",
          7933 => x"81",
          7934 => x"b6",
          7935 => x"78",
          7936 => x"3f",
          7937 => x"08",
          7938 => x"98",
          7939 => x"38",
          7940 => x"52",
          7941 => x"ff",
          7942 => x"78",
          7943 => x"b4",
          7944 => x"54",
          7945 => x"15",
          7946 => x"b2",
          7947 => x"ca",
          7948 => x"b6",
          7949 => x"53",
          7950 => x"53",
          7951 => x"3f",
          7952 => x"b4",
          7953 => x"d4",
          7954 => x"b6",
          7955 => x"54",
          7956 => x"d5",
          7957 => x"53",
          7958 => x"11",
          7959 => x"d7",
          7960 => x"81",
          7961 => x"34",
          7962 => x"a4",
          7963 => x"98",
          7964 => x"b6",
          7965 => x"38",
          7966 => x"0a",
          7967 => x"05",
          7968 => x"d0",
          7969 => x"64",
          7970 => x"c9",
          7971 => x"54",
          7972 => x"15",
          7973 => x"81",
          7974 => x"34",
          7975 => x"b8",
          7976 => x"b6",
          7977 => x"8b",
          7978 => x"75",
          7979 => x"ff",
          7980 => x"73",
          7981 => x"0c",
          7982 => x"04",
          7983 => x"a9",
          7984 => x"51",
          7985 => x"82",
          7986 => x"ff",
          7987 => x"a9",
          7988 => x"ee",
          7989 => x"98",
          7990 => x"b6",
          7991 => x"d3",
          7992 => x"a9",
          7993 => x"9d",
          7994 => x"58",
          7995 => x"82",
          7996 => x"55",
          7997 => x"08",
          7998 => x"02",
          7999 => x"33",
          8000 => x"54",
          8001 => x"82",
          8002 => x"53",
          8003 => x"52",
          8004 => x"88",
          8005 => x"b4",
          8006 => x"53",
          8007 => x"3d",
          8008 => x"ff",
          8009 => x"aa",
          8010 => x"73",
          8011 => x"3f",
          8012 => x"08",
          8013 => x"98",
          8014 => x"63",
          8015 => x"81",
          8016 => x"65",
          8017 => x"2e",
          8018 => x"55",
          8019 => x"82",
          8020 => x"84",
          8021 => x"06",
          8022 => x"73",
          8023 => x"3f",
          8024 => x"08",
          8025 => x"98",
          8026 => x"38",
          8027 => x"53",
          8028 => x"95",
          8029 => x"16",
          8030 => x"87",
          8031 => x"05",
          8032 => x"34",
          8033 => x"70",
          8034 => x"81",
          8035 => x"55",
          8036 => x"74",
          8037 => x"73",
          8038 => x"78",
          8039 => x"83",
          8040 => x"16",
          8041 => x"2a",
          8042 => x"51",
          8043 => x"80",
          8044 => x"38",
          8045 => x"80",
          8046 => x"52",
          8047 => x"be",
          8048 => x"98",
          8049 => x"51",
          8050 => x"3f",
          8051 => x"b6",
          8052 => x"2e",
          8053 => x"82",
          8054 => x"52",
          8055 => x"b5",
          8056 => x"b6",
          8057 => x"80",
          8058 => x"58",
          8059 => x"98",
          8060 => x"38",
          8061 => x"54",
          8062 => x"09",
          8063 => x"38",
          8064 => x"52",
          8065 => x"af",
          8066 => x"81",
          8067 => x"34",
          8068 => x"b6",
          8069 => x"38",
          8070 => x"ca",
          8071 => x"98",
          8072 => x"b6",
          8073 => x"38",
          8074 => x"b5",
          8075 => x"b6",
          8076 => x"74",
          8077 => x"0c",
          8078 => x"04",
          8079 => x"02",
          8080 => x"33",
          8081 => x"80",
          8082 => x"57",
          8083 => x"95",
          8084 => x"52",
          8085 => x"d2",
          8086 => x"b6",
          8087 => x"82",
          8088 => x"80",
          8089 => x"5a",
          8090 => x"3d",
          8091 => x"c9",
          8092 => x"b6",
          8093 => x"82",
          8094 => x"b8",
          8095 => x"cf",
          8096 => x"a0",
          8097 => x"55",
          8098 => x"75",
          8099 => x"71",
          8100 => x"33",
          8101 => x"74",
          8102 => x"57",
          8103 => x"8b",
          8104 => x"54",
          8105 => x"15",
          8106 => x"ff",
          8107 => x"82",
          8108 => x"55",
          8109 => x"98",
          8110 => x"0d",
          8111 => x"0d",
          8112 => x"53",
          8113 => x"05",
          8114 => x"51",
          8115 => x"82",
          8116 => x"55",
          8117 => x"08",
          8118 => x"76",
          8119 => x"93",
          8120 => x"51",
          8121 => x"82",
          8122 => x"55",
          8123 => x"08",
          8124 => x"80",
          8125 => x"81",
          8126 => x"86",
          8127 => x"38",
          8128 => x"86",
          8129 => x"90",
          8130 => x"54",
          8131 => x"ff",
          8132 => x"76",
          8133 => x"83",
          8134 => x"51",
          8135 => x"3f",
          8136 => x"08",
          8137 => x"b6",
          8138 => x"3d",
          8139 => x"3d",
          8140 => x"5c",
          8141 => x"98",
          8142 => x"52",
          8143 => x"d1",
          8144 => x"b6",
          8145 => x"b6",
          8146 => x"70",
          8147 => x"08",
          8148 => x"51",
          8149 => x"80",
          8150 => x"38",
          8151 => x"06",
          8152 => x"80",
          8153 => x"38",
          8154 => x"5f",
          8155 => x"3d",
          8156 => x"ff",
          8157 => x"82",
          8158 => x"57",
          8159 => x"08",
          8160 => x"74",
          8161 => x"c3",
          8162 => x"b6",
          8163 => x"82",
          8164 => x"bf",
          8165 => x"98",
          8166 => x"98",
          8167 => x"59",
          8168 => x"81",
          8169 => x"56",
          8170 => x"33",
          8171 => x"16",
          8172 => x"27",
          8173 => x"56",
          8174 => x"80",
          8175 => x"80",
          8176 => x"ff",
          8177 => x"70",
          8178 => x"56",
          8179 => x"e8",
          8180 => x"76",
          8181 => x"81",
          8182 => x"80",
          8183 => x"57",
          8184 => x"78",
          8185 => x"51",
          8186 => x"2e",
          8187 => x"73",
          8188 => x"38",
          8189 => x"08",
          8190 => x"b1",
          8191 => x"b6",
          8192 => x"82",
          8193 => x"a7",
          8194 => x"33",
          8195 => x"c3",
          8196 => x"2e",
          8197 => x"e4",
          8198 => x"2e",
          8199 => x"56",
          8200 => x"05",
          8201 => x"e3",
          8202 => x"98",
          8203 => x"76",
          8204 => x"0c",
          8205 => x"04",
          8206 => x"82",
          8207 => x"ff",
          8208 => x"9d",
          8209 => x"fa",
          8210 => x"98",
          8211 => x"98",
          8212 => x"82",
          8213 => x"83",
          8214 => x"53",
          8215 => x"3d",
          8216 => x"ff",
          8217 => x"73",
          8218 => x"70",
          8219 => x"52",
          8220 => x"9f",
          8221 => x"bc",
          8222 => x"74",
          8223 => x"6d",
          8224 => x"70",
          8225 => x"af",
          8226 => x"b6",
          8227 => x"2e",
          8228 => x"70",
          8229 => x"57",
          8230 => x"fd",
          8231 => x"98",
          8232 => x"8d",
          8233 => x"2b",
          8234 => x"81",
          8235 => x"86",
          8236 => x"98",
          8237 => x"9f",
          8238 => x"ff",
          8239 => x"54",
          8240 => x"8a",
          8241 => x"70",
          8242 => x"06",
          8243 => x"ff",
          8244 => x"38",
          8245 => x"15",
          8246 => x"80",
          8247 => x"74",
          8248 => x"e0",
          8249 => x"89",
          8250 => x"98",
          8251 => x"81",
          8252 => x"88",
          8253 => x"26",
          8254 => x"39",
          8255 => x"86",
          8256 => x"81",
          8257 => x"ff",
          8258 => x"38",
          8259 => x"54",
          8260 => x"81",
          8261 => x"81",
          8262 => x"78",
          8263 => x"5a",
          8264 => x"6d",
          8265 => x"81",
          8266 => x"57",
          8267 => x"9f",
          8268 => x"38",
          8269 => x"54",
          8270 => x"81",
          8271 => x"b1",
          8272 => x"2e",
          8273 => x"a7",
          8274 => x"15",
          8275 => x"54",
          8276 => x"09",
          8277 => x"38",
          8278 => x"76",
          8279 => x"41",
          8280 => x"52",
          8281 => x"52",
          8282 => x"b3",
          8283 => x"98",
          8284 => x"b6",
          8285 => x"f7",
          8286 => x"74",
          8287 => x"e5",
          8288 => x"98",
          8289 => x"b6",
          8290 => x"38",
          8291 => x"38",
          8292 => x"74",
          8293 => x"39",
          8294 => x"08",
          8295 => x"81",
          8296 => x"38",
          8297 => x"74",
          8298 => x"38",
          8299 => x"51",
          8300 => x"3f",
          8301 => x"08",
          8302 => x"98",
          8303 => x"a0",
          8304 => x"98",
          8305 => x"51",
          8306 => x"3f",
          8307 => x"0b",
          8308 => x"8b",
          8309 => x"67",
          8310 => x"a7",
          8311 => x"81",
          8312 => x"34",
          8313 => x"ad",
          8314 => x"b6",
          8315 => x"73",
          8316 => x"b6",
          8317 => x"3d",
          8318 => x"3d",
          8319 => x"02",
          8320 => x"cb",
          8321 => x"3d",
          8322 => x"72",
          8323 => x"5a",
          8324 => x"82",
          8325 => x"58",
          8326 => x"08",
          8327 => x"91",
          8328 => x"77",
          8329 => x"7c",
          8330 => x"38",
          8331 => x"59",
          8332 => x"90",
          8333 => x"81",
          8334 => x"06",
          8335 => x"73",
          8336 => x"54",
          8337 => x"82",
          8338 => x"39",
          8339 => x"8b",
          8340 => x"11",
          8341 => x"2b",
          8342 => x"54",
          8343 => x"fe",
          8344 => x"ff",
          8345 => x"70",
          8346 => x"07",
          8347 => x"b6",
          8348 => x"8c",
          8349 => x"40",
          8350 => x"55",
          8351 => x"88",
          8352 => x"08",
          8353 => x"38",
          8354 => x"77",
          8355 => x"56",
          8356 => x"51",
          8357 => x"3f",
          8358 => x"55",
          8359 => x"08",
          8360 => x"38",
          8361 => x"b6",
          8362 => x"2e",
          8363 => x"82",
          8364 => x"ff",
          8365 => x"38",
          8366 => x"08",
          8367 => x"16",
          8368 => x"2e",
          8369 => x"87",
          8370 => x"74",
          8371 => x"74",
          8372 => x"81",
          8373 => x"38",
          8374 => x"ff",
          8375 => x"2e",
          8376 => x"7b",
          8377 => x"80",
          8378 => x"81",
          8379 => x"81",
          8380 => x"06",
          8381 => x"56",
          8382 => x"52",
          8383 => x"af",
          8384 => x"b6",
          8385 => x"82",
          8386 => x"80",
          8387 => x"81",
          8388 => x"56",
          8389 => x"d3",
          8390 => x"ff",
          8391 => x"7c",
          8392 => x"55",
          8393 => x"b3",
          8394 => x"1b",
          8395 => x"1b",
          8396 => x"33",
          8397 => x"54",
          8398 => x"34",
          8399 => x"fe",
          8400 => x"08",
          8401 => x"74",
          8402 => x"75",
          8403 => x"16",
          8404 => x"33",
          8405 => x"73",
          8406 => x"77",
          8407 => x"b6",
          8408 => x"3d",
          8409 => x"3d",
          8410 => x"02",
          8411 => x"eb",
          8412 => x"3d",
          8413 => x"59",
          8414 => x"8b",
          8415 => x"82",
          8416 => x"24",
          8417 => x"82",
          8418 => x"84",
          8419 => x"d0",
          8420 => x"51",
          8421 => x"2e",
          8422 => x"75",
          8423 => x"98",
          8424 => x"06",
          8425 => x"7e",
          8426 => x"d0",
          8427 => x"98",
          8428 => x"06",
          8429 => x"56",
          8430 => x"74",
          8431 => x"76",
          8432 => x"81",
          8433 => x"8a",
          8434 => x"b2",
          8435 => x"fc",
          8436 => x"52",
          8437 => x"a4",
          8438 => x"b6",
          8439 => x"38",
          8440 => x"80",
          8441 => x"74",
          8442 => x"26",
          8443 => x"15",
          8444 => x"74",
          8445 => x"38",
          8446 => x"80",
          8447 => x"84",
          8448 => x"92",
          8449 => x"80",
          8450 => x"38",
          8451 => x"06",
          8452 => x"2e",
          8453 => x"56",
          8454 => x"78",
          8455 => x"89",
          8456 => x"2b",
          8457 => x"43",
          8458 => x"38",
          8459 => x"30",
          8460 => x"77",
          8461 => x"91",
          8462 => x"c2",
          8463 => x"f8",
          8464 => x"52",
          8465 => x"a4",
          8466 => x"56",
          8467 => x"08",
          8468 => x"77",
          8469 => x"77",
          8470 => x"98",
          8471 => x"45",
          8472 => x"bf",
          8473 => x"8e",
          8474 => x"26",
          8475 => x"74",
          8476 => x"48",
          8477 => x"75",
          8478 => x"38",
          8479 => x"81",
          8480 => x"fa",
          8481 => x"2a",
          8482 => x"56",
          8483 => x"2e",
          8484 => x"87",
          8485 => x"82",
          8486 => x"38",
          8487 => x"55",
          8488 => x"83",
          8489 => x"81",
          8490 => x"56",
          8491 => x"80",
          8492 => x"38",
          8493 => x"83",
          8494 => x"06",
          8495 => x"78",
          8496 => x"91",
          8497 => x"0b",
          8498 => x"22",
          8499 => x"80",
          8500 => x"74",
          8501 => x"38",
          8502 => x"56",
          8503 => x"17",
          8504 => x"57",
          8505 => x"2e",
          8506 => x"75",
          8507 => x"79",
          8508 => x"fe",
          8509 => x"82",
          8510 => x"84",
          8511 => x"05",
          8512 => x"5e",
          8513 => x"80",
          8514 => x"98",
          8515 => x"8a",
          8516 => x"fd",
          8517 => x"75",
          8518 => x"38",
          8519 => x"78",
          8520 => x"8c",
          8521 => x"0b",
          8522 => x"22",
          8523 => x"80",
          8524 => x"74",
          8525 => x"38",
          8526 => x"56",
          8527 => x"17",
          8528 => x"57",
          8529 => x"2e",
          8530 => x"75",
          8531 => x"79",
          8532 => x"fe",
          8533 => x"82",
          8534 => x"10",
          8535 => x"82",
          8536 => x"9f",
          8537 => x"38",
          8538 => x"b6",
          8539 => x"82",
          8540 => x"05",
          8541 => x"2a",
          8542 => x"56",
          8543 => x"17",
          8544 => x"81",
          8545 => x"60",
          8546 => x"65",
          8547 => x"12",
          8548 => x"30",
          8549 => x"74",
          8550 => x"59",
          8551 => x"7d",
          8552 => x"81",
          8553 => x"76",
          8554 => x"41",
          8555 => x"76",
          8556 => x"90",
          8557 => x"62",
          8558 => x"51",
          8559 => x"26",
          8560 => x"75",
          8561 => x"31",
          8562 => x"65",
          8563 => x"fe",
          8564 => x"82",
          8565 => x"58",
          8566 => x"09",
          8567 => x"38",
          8568 => x"08",
          8569 => x"26",
          8570 => x"78",
          8571 => x"79",
          8572 => x"78",
          8573 => x"86",
          8574 => x"82",
          8575 => x"06",
          8576 => x"83",
          8577 => x"82",
          8578 => x"27",
          8579 => x"8f",
          8580 => x"55",
          8581 => x"26",
          8582 => x"59",
          8583 => x"62",
          8584 => x"74",
          8585 => x"38",
          8586 => x"88",
          8587 => x"98",
          8588 => x"26",
          8589 => x"86",
          8590 => x"1a",
          8591 => x"79",
          8592 => x"38",
          8593 => x"80",
          8594 => x"2e",
          8595 => x"83",
          8596 => x"9f",
          8597 => x"8b",
          8598 => x"06",
          8599 => x"74",
          8600 => x"84",
          8601 => x"52",
          8602 => x"a2",
          8603 => x"53",
          8604 => x"52",
          8605 => x"a2",
          8606 => x"80",
          8607 => x"51",
          8608 => x"3f",
          8609 => x"34",
          8610 => x"ff",
          8611 => x"1b",
          8612 => x"a2",
          8613 => x"90",
          8614 => x"83",
          8615 => x"70",
          8616 => x"80",
          8617 => x"55",
          8618 => x"ff",
          8619 => x"66",
          8620 => x"ff",
          8621 => x"38",
          8622 => x"ff",
          8623 => x"1b",
          8624 => x"f2",
          8625 => x"74",
          8626 => x"51",
          8627 => x"3f",
          8628 => x"1c",
          8629 => x"98",
          8630 => x"a0",
          8631 => x"ff",
          8632 => x"51",
          8633 => x"3f",
          8634 => x"1b",
          8635 => x"e4",
          8636 => x"2e",
          8637 => x"80",
          8638 => x"88",
          8639 => x"80",
          8640 => x"ff",
          8641 => x"7c",
          8642 => x"51",
          8643 => x"3f",
          8644 => x"1b",
          8645 => x"bc",
          8646 => x"b0",
          8647 => x"a0",
          8648 => x"52",
          8649 => x"ff",
          8650 => x"ff",
          8651 => x"c0",
          8652 => x"0b",
          8653 => x"34",
          8654 => x"af",
          8655 => x"c7",
          8656 => x"39",
          8657 => x"0a",
          8658 => x"51",
          8659 => x"3f",
          8660 => x"ff",
          8661 => x"1b",
          8662 => x"da",
          8663 => x"0b",
          8664 => x"a9",
          8665 => x"34",
          8666 => x"af",
          8667 => x"1b",
          8668 => x"8f",
          8669 => x"d5",
          8670 => x"1b",
          8671 => x"ff",
          8672 => x"81",
          8673 => x"7a",
          8674 => x"ff",
          8675 => x"81",
          8676 => x"98",
          8677 => x"38",
          8678 => x"09",
          8679 => x"ee",
          8680 => x"60",
          8681 => x"7a",
          8682 => x"ff",
          8683 => x"84",
          8684 => x"52",
          8685 => x"9f",
          8686 => x"8b",
          8687 => x"52",
          8688 => x"9f",
          8689 => x"8a",
          8690 => x"52",
          8691 => x"51",
          8692 => x"3f",
          8693 => x"83",
          8694 => x"ff",
          8695 => x"82",
          8696 => x"1b",
          8697 => x"ec",
          8698 => x"d5",
          8699 => x"ff",
          8700 => x"75",
          8701 => x"05",
          8702 => x"7e",
          8703 => x"e5",
          8704 => x"60",
          8705 => x"52",
          8706 => x"9a",
          8707 => x"53",
          8708 => x"51",
          8709 => x"3f",
          8710 => x"58",
          8711 => x"09",
          8712 => x"38",
          8713 => x"51",
          8714 => x"3f",
          8715 => x"1b",
          8716 => x"a0",
          8717 => x"52",
          8718 => x"91",
          8719 => x"ff",
          8720 => x"81",
          8721 => x"f8",
          8722 => x"7a",
          8723 => x"84",
          8724 => x"61",
          8725 => x"26",
          8726 => x"57",
          8727 => x"53",
          8728 => x"51",
          8729 => x"3f",
          8730 => x"08",
          8731 => x"84",
          8732 => x"b6",
          8733 => x"7a",
          8734 => x"aa",
          8735 => x"75",
          8736 => x"56",
          8737 => x"81",
          8738 => x"80",
          8739 => x"38",
          8740 => x"83",
          8741 => x"63",
          8742 => x"74",
          8743 => x"38",
          8744 => x"54",
          8745 => x"52",
          8746 => x"99",
          8747 => x"b6",
          8748 => x"c1",
          8749 => x"75",
          8750 => x"56",
          8751 => x"8c",
          8752 => x"2e",
          8753 => x"56",
          8754 => x"ff",
          8755 => x"84",
          8756 => x"2e",
          8757 => x"56",
          8758 => x"58",
          8759 => x"38",
          8760 => x"77",
          8761 => x"ff",
          8762 => x"82",
          8763 => x"78",
          8764 => x"c2",
          8765 => x"1b",
          8766 => x"34",
          8767 => x"16",
          8768 => x"82",
          8769 => x"83",
          8770 => x"84",
          8771 => x"67",
          8772 => x"fd",
          8773 => x"51",
          8774 => x"3f",
          8775 => x"16",
          8776 => x"98",
          8777 => x"bf",
          8778 => x"86",
          8779 => x"b6",
          8780 => x"16",
          8781 => x"83",
          8782 => x"ff",
          8783 => x"66",
          8784 => x"1b",
          8785 => x"8c",
          8786 => x"77",
          8787 => x"7e",
          8788 => x"91",
          8789 => x"82",
          8790 => x"a2",
          8791 => x"80",
          8792 => x"ff",
          8793 => x"81",
          8794 => x"98",
          8795 => x"89",
          8796 => x"8a",
          8797 => x"86",
          8798 => x"98",
          8799 => x"82",
          8800 => x"99",
          8801 => x"f5",
          8802 => x"60",
          8803 => x"79",
          8804 => x"5a",
          8805 => x"78",
          8806 => x"8d",
          8807 => x"55",
          8808 => x"fc",
          8809 => x"51",
          8810 => x"7a",
          8811 => x"81",
          8812 => x"8c",
          8813 => x"74",
          8814 => x"38",
          8815 => x"81",
          8816 => x"81",
          8817 => x"8a",
          8818 => x"06",
          8819 => x"76",
          8820 => x"76",
          8821 => x"55",
          8822 => x"98",
          8823 => x"0d",
          8824 => x"0d",
          8825 => x"05",
          8826 => x"59",
          8827 => x"2e",
          8828 => x"87",
          8829 => x"76",
          8830 => x"84",
          8831 => x"80",
          8832 => x"38",
          8833 => x"77",
          8834 => x"56",
          8835 => x"34",
          8836 => x"bb",
          8837 => x"38",
          8838 => x"05",
          8839 => x"8c",
          8840 => x"08",
          8841 => x"3f",
          8842 => x"70",
          8843 => x"07",
          8844 => x"30",
          8845 => x"56",
          8846 => x"0c",
          8847 => x"18",
          8848 => x"0d",
          8849 => x"0d",
          8850 => x"08",
          8851 => x"75",
          8852 => x"89",
          8853 => x"54",
          8854 => x"16",
          8855 => x"51",
          8856 => x"82",
          8857 => x"91",
          8858 => x"08",
          8859 => x"81",
          8860 => x"88",
          8861 => x"83",
          8862 => x"74",
          8863 => x"0c",
          8864 => x"04",
          8865 => x"75",
          8866 => x"53",
          8867 => x"51",
          8868 => x"3f",
          8869 => x"85",
          8870 => x"ea",
          8871 => x"80",
          8872 => x"6a",
          8873 => x"70",
          8874 => x"d8",
          8875 => x"72",
          8876 => x"3f",
          8877 => x"8d",
          8878 => x"0d",
          8879 => x"00",
          8880 => x"ff",
          8881 => x"ff",
          8882 => x"ff",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"64",
          9020 => x"74",
          9021 => x"64",
          9022 => x"74",
          9023 => x"66",
          9024 => x"74",
          9025 => x"66",
          9026 => x"64",
          9027 => x"66",
          9028 => x"63",
          9029 => x"6d",
          9030 => x"61",
          9031 => x"6d",
          9032 => x"79",
          9033 => x"6d",
          9034 => x"66",
          9035 => x"6d",
          9036 => x"70",
          9037 => x"6d",
          9038 => x"6d",
          9039 => x"6d",
          9040 => x"68",
          9041 => x"68",
          9042 => x"68",
          9043 => x"68",
          9044 => x"63",
          9045 => x"00",
          9046 => x"6a",
          9047 => x"72",
          9048 => x"61",
          9049 => x"72",
          9050 => x"74",
          9051 => x"69",
          9052 => x"00",
          9053 => x"74",
          9054 => x"00",
          9055 => x"74",
          9056 => x"69",
          9057 => x"6d",
          9058 => x"69",
          9059 => x"6b",
          9060 => x"00",
          9061 => x"65",
          9062 => x"44",
          9063 => x"20",
          9064 => x"6f",
          9065 => x"49",
          9066 => x"72",
          9067 => x"20",
          9068 => x"6f",
          9069 => x"44",
          9070 => x"20",
          9071 => x"20",
          9072 => x"64",
          9073 => x"4e",
          9074 => x"69",
          9075 => x"66",
          9076 => x"64",
          9077 => x"4e",
          9078 => x"61",
          9079 => x"66",
          9080 => x"64",
          9081 => x"49",
          9082 => x"6c",
          9083 => x"66",
          9084 => x"6e",
          9085 => x"2e",
          9086 => x"41",
          9087 => x"73",
          9088 => x"65",
          9089 => x"64",
          9090 => x"46",
          9091 => x"20",
          9092 => x"65",
          9093 => x"20",
          9094 => x"73",
          9095 => x"00",
          9096 => x"46",
          9097 => x"20",
          9098 => x"64",
          9099 => x"69",
          9100 => x"6c",
          9101 => x"00",
          9102 => x"53",
          9103 => x"73",
          9104 => x"69",
          9105 => x"70",
          9106 => x"65",
          9107 => x"64",
          9108 => x"44",
          9109 => x"65",
          9110 => x"6d",
          9111 => x"20",
          9112 => x"69",
          9113 => x"6c",
          9114 => x"00",
          9115 => x"44",
          9116 => x"20",
          9117 => x"20",
          9118 => x"62",
          9119 => x"2e",
          9120 => x"4e",
          9121 => x"6f",
          9122 => x"74",
          9123 => x"65",
          9124 => x"6c",
          9125 => x"73",
          9126 => x"20",
          9127 => x"6e",
          9128 => x"6e",
          9129 => x"73",
          9130 => x"46",
          9131 => x"61",
          9132 => x"62",
          9133 => x"65",
          9134 => x"54",
          9135 => x"6f",
          9136 => x"20",
          9137 => x"72",
          9138 => x"6f",
          9139 => x"61",
          9140 => x"6c",
          9141 => x"2e",
          9142 => x"46",
          9143 => x"20",
          9144 => x"6c",
          9145 => x"65",
          9146 => x"49",
          9147 => x"66",
          9148 => x"69",
          9149 => x"20",
          9150 => x"6f",
          9151 => x"00",
          9152 => x"54",
          9153 => x"6d",
          9154 => x"20",
          9155 => x"6e",
          9156 => x"6c",
          9157 => x"00",
          9158 => x"50",
          9159 => x"6d",
          9160 => x"72",
          9161 => x"6e",
          9162 => x"72",
          9163 => x"2e",
          9164 => x"53",
          9165 => x"65",
          9166 => x"00",
          9167 => x"55",
          9168 => x"6f",
          9169 => x"65",
          9170 => x"72",
          9171 => x"0a",
          9172 => x"20",
          9173 => x"65",
          9174 => x"73",
          9175 => x"20",
          9176 => x"20",
          9177 => x"65",
          9178 => x"65",
          9179 => x"00",
          9180 => x"72",
          9181 => x"00",
          9182 => x"30",
          9183 => x"38",
          9184 => x"20",
          9185 => x"30",
          9186 => x"2c",
          9187 => x"25",
          9188 => x"78",
          9189 => x"49",
          9190 => x"25",
          9191 => x"78",
          9192 => x"38",
          9193 => x"25",
          9194 => x"78",
          9195 => x"25",
          9196 => x"58",
          9197 => x"3a",
          9198 => x"25",
          9199 => x"00",
          9200 => x"20",
          9201 => x"20",
          9202 => x"00",
          9203 => x"25",
          9204 => x"00",
          9205 => x"20",
          9206 => x"20",
          9207 => x"7c",
          9208 => x"7a",
          9209 => x"0a",
          9210 => x"25",
          9211 => x"00",
          9212 => x"30",
          9213 => x"35",
          9214 => x"32",
          9215 => x"76",
          9216 => x"32",
          9217 => x"20",
          9218 => x"2c",
          9219 => x"76",
          9220 => x"32",
          9221 => x"25",
          9222 => x"73",
          9223 => x"0a",
          9224 => x"5a",
          9225 => x"49",
          9226 => x"72",
          9227 => x"74",
          9228 => x"6e",
          9229 => x"72",
          9230 => x"54",
          9231 => x"72",
          9232 => x"74",
          9233 => x"75",
          9234 => x"50",
          9235 => x"69",
          9236 => x"72",
          9237 => x"74",
          9238 => x"49",
          9239 => x"4c",
          9240 => x"20",
          9241 => x"65",
          9242 => x"70",
          9243 => x"49",
          9244 => x"4c",
          9245 => x"20",
          9246 => x"65",
          9247 => x"70",
          9248 => x"55",
          9249 => x"30",
          9250 => x"20",
          9251 => x"65",
          9252 => x"70",
          9253 => x"55",
          9254 => x"30",
          9255 => x"20",
          9256 => x"65",
          9257 => x"70",
          9258 => x"55",
          9259 => x"31",
          9260 => x"20",
          9261 => x"65",
          9262 => x"70",
          9263 => x"55",
          9264 => x"31",
          9265 => x"20",
          9266 => x"65",
          9267 => x"70",
          9268 => x"53",
          9269 => x"69",
          9270 => x"75",
          9271 => x"69",
          9272 => x"2e",
          9273 => x"45",
          9274 => x"6c",
          9275 => x"20",
          9276 => x"65",
          9277 => x"2e",
          9278 => x"61",
          9279 => x"65",
          9280 => x"2e",
          9281 => x"00",
          9282 => x"7a",
          9283 => x"68",
          9284 => x"30",
          9285 => x"46",
          9286 => x"65",
          9287 => x"6f",
          9288 => x"69",
          9289 => x"6c",
          9290 => x"20",
          9291 => x"63",
          9292 => x"20",
          9293 => x"70",
          9294 => x"73",
          9295 => x"6e",
          9296 => x"6d",
          9297 => x"61",
          9298 => x"2e",
          9299 => x"2a",
          9300 => x"43",
          9301 => x"72",
          9302 => x"2e",
          9303 => x"00",
          9304 => x"43",
          9305 => x"69",
          9306 => x"2e",
          9307 => x"43",
          9308 => x"61",
          9309 => x"67",
          9310 => x"00",
          9311 => x"25",
          9312 => x"78",
          9313 => x"38",
          9314 => x"3e",
          9315 => x"6c",
          9316 => x"30",
          9317 => x"0a",
          9318 => x"44",
          9319 => x"20",
          9320 => x"6f",
          9321 => x"0a",
          9322 => x"70",
          9323 => x"65",
          9324 => x"25",
          9325 => x"58",
          9326 => x"32",
          9327 => x"3f",
          9328 => x"25",
          9329 => x"58",
          9330 => x"34",
          9331 => x"25",
          9332 => x"58",
          9333 => x"38",
          9334 => x"00",
          9335 => x"45",
          9336 => x"75",
          9337 => x"67",
          9338 => x"64",
          9339 => x"20",
          9340 => x"6c",
          9341 => x"2e",
          9342 => x"43",
          9343 => x"69",
          9344 => x"63",
          9345 => x"20",
          9346 => x"30",
          9347 => x"20",
          9348 => x"0a",
          9349 => x"43",
          9350 => x"20",
          9351 => x"75",
          9352 => x"64",
          9353 => x"64",
          9354 => x"25",
          9355 => x"0a",
          9356 => x"52",
          9357 => x"61",
          9358 => x"6e",
          9359 => x"70",
          9360 => x"63",
          9361 => x"6f",
          9362 => x"2e",
          9363 => x"43",
          9364 => x"20",
          9365 => x"6f",
          9366 => x"6e",
          9367 => x"2e",
          9368 => x"5a",
          9369 => x"62",
          9370 => x"25",
          9371 => x"25",
          9372 => x"73",
          9373 => x"00",
          9374 => x"25",
          9375 => x"25",
          9376 => x"73",
          9377 => x"25",
          9378 => x"25",
          9379 => x"42",
          9380 => x"63",
          9381 => x"61",
          9382 => x"00",
          9383 => x"52",
          9384 => x"69",
          9385 => x"2e",
          9386 => x"45",
          9387 => x"6c",
          9388 => x"20",
          9389 => x"65",
          9390 => x"70",
          9391 => x"2e",
          9392 => x"25",
          9393 => x"64",
          9394 => x"20",
          9395 => x"25",
          9396 => x"64",
          9397 => x"25",
          9398 => x"53",
          9399 => x"43",
          9400 => x"69",
          9401 => x"61",
          9402 => x"6e",
          9403 => x"20",
          9404 => x"6f",
          9405 => x"6f",
          9406 => x"6f",
          9407 => x"67",
          9408 => x"3a",
          9409 => x"76",
          9410 => x"73",
          9411 => x"70",
          9412 => x"65",
          9413 => x"64",
          9414 => x"20",
          9415 => x"57",
          9416 => x"44",
          9417 => x"20",
          9418 => x"30",
          9419 => x"25",
          9420 => x"29",
          9421 => x"20",
          9422 => x"53",
          9423 => x"4d",
          9424 => x"20",
          9425 => x"30",
          9426 => x"25",
          9427 => x"29",
          9428 => x"20",
          9429 => x"49",
          9430 => x"20",
          9431 => x"4d",
          9432 => x"30",
          9433 => x"25",
          9434 => x"29",
          9435 => x"20",
          9436 => x"42",
          9437 => x"20",
          9438 => x"20",
          9439 => x"30",
          9440 => x"25",
          9441 => x"29",
          9442 => x"20",
          9443 => x"52",
          9444 => x"20",
          9445 => x"20",
          9446 => x"30",
          9447 => x"25",
          9448 => x"29",
          9449 => x"20",
          9450 => x"53",
          9451 => x"41",
          9452 => x"20",
          9453 => x"65",
          9454 => x"65",
          9455 => x"25",
          9456 => x"29",
          9457 => x"20",
          9458 => x"54",
          9459 => x"52",
          9460 => x"20",
          9461 => x"69",
          9462 => x"73",
          9463 => x"25",
          9464 => x"29",
          9465 => x"20",
          9466 => x"49",
          9467 => x"20",
          9468 => x"4c",
          9469 => x"68",
          9470 => x"65",
          9471 => x"25",
          9472 => x"29",
          9473 => x"20",
          9474 => x"57",
          9475 => x"42",
          9476 => x"20",
          9477 => x"00",
          9478 => x"20",
          9479 => x"57",
          9480 => x"32",
          9481 => x"20",
          9482 => x"49",
          9483 => x"4c",
          9484 => x"20",
          9485 => x"50",
          9486 => x"20",
          9487 => x"53",
          9488 => x"41",
          9489 => x"65",
          9490 => x"73",
          9491 => x"20",
          9492 => x"43",
          9493 => x"52",
          9494 => x"74",
          9495 => x"63",
          9496 => x"20",
          9497 => x"72",
          9498 => x"20",
          9499 => x"30",
          9500 => x"00",
          9501 => x"20",
          9502 => x"43",
          9503 => x"4d",
          9504 => x"72",
          9505 => x"74",
          9506 => x"20",
          9507 => x"72",
          9508 => x"20",
          9509 => x"30",
          9510 => x"00",
          9511 => x"20",
          9512 => x"53",
          9513 => x"6b",
          9514 => x"61",
          9515 => x"41",
          9516 => x"65",
          9517 => x"20",
          9518 => x"20",
          9519 => x"30",
          9520 => x"00",
          9521 => x"4d",
          9522 => x"3a",
          9523 => x"20",
          9524 => x"5a",
          9525 => x"49",
          9526 => x"20",
          9527 => x"20",
          9528 => x"20",
          9529 => x"20",
          9530 => x"20",
          9531 => x"30",
          9532 => x"00",
          9533 => x"20",
          9534 => x"53",
          9535 => x"65",
          9536 => x"6c",
          9537 => x"20",
          9538 => x"71",
          9539 => x"20",
          9540 => x"20",
          9541 => x"64",
          9542 => x"34",
          9543 => x"7a",
          9544 => x"20",
          9545 => x"53",
          9546 => x"4d",
          9547 => x"6f",
          9548 => x"46",
          9549 => x"20",
          9550 => x"20",
          9551 => x"20",
          9552 => x"64",
          9553 => x"34",
          9554 => x"7a",
          9555 => x"20",
          9556 => x"57",
          9557 => x"62",
          9558 => x"20",
          9559 => x"41",
          9560 => x"6c",
          9561 => x"20",
          9562 => x"71",
          9563 => x"64",
          9564 => x"34",
          9565 => x"7a",
          9566 => x"53",
          9567 => x"6c",
          9568 => x"4d",
          9569 => x"75",
          9570 => x"46",
          9571 => x"00",
          9572 => x"45",
          9573 => x"45",
          9574 => x"00",
          9575 => x"55",
          9576 => x"6f",
          9577 => x"00",
          9578 => x"01",
          9579 => x"00",
          9580 => x"00",
          9581 => x"01",
          9582 => x"00",
          9583 => x"00",
          9584 => x"01",
          9585 => x"00",
          9586 => x"00",
          9587 => x"01",
          9588 => x"00",
          9589 => x"00",
          9590 => x"01",
          9591 => x"00",
          9592 => x"00",
          9593 => x"01",
          9594 => x"00",
          9595 => x"00",
          9596 => x"01",
          9597 => x"00",
          9598 => x"00",
          9599 => x"01",
          9600 => x"00",
          9601 => x"00",
          9602 => x"01",
          9603 => x"00",
          9604 => x"00",
          9605 => x"01",
          9606 => x"00",
          9607 => x"00",
          9608 => x"01",
          9609 => x"00",
          9610 => x"00",
          9611 => x"04",
          9612 => x"00",
          9613 => x"00",
          9614 => x"04",
          9615 => x"00",
          9616 => x"00",
          9617 => x"04",
          9618 => x"00",
          9619 => x"00",
          9620 => x"03",
          9621 => x"00",
          9622 => x"00",
          9623 => x"04",
          9624 => x"00",
          9625 => x"00",
          9626 => x"04",
          9627 => x"00",
          9628 => x"00",
          9629 => x"04",
          9630 => x"00",
          9631 => x"00",
          9632 => x"03",
          9633 => x"00",
          9634 => x"00",
          9635 => x"03",
          9636 => x"00",
          9637 => x"00",
          9638 => x"03",
          9639 => x"00",
          9640 => x"00",
          9641 => x"03",
          9642 => x"00",
          9643 => x"1b",
          9644 => x"1b",
          9645 => x"1b",
          9646 => x"1b",
          9647 => x"1b",
          9648 => x"1b",
          9649 => x"1b",
          9650 => x"1b",
          9651 => x"1b",
          9652 => x"1b",
          9653 => x"1b",
          9654 => x"10",
          9655 => x"0e",
          9656 => x"0d",
          9657 => x"0b",
          9658 => x"08",
          9659 => x"06",
          9660 => x"05",
          9661 => x"04",
          9662 => x"03",
          9663 => x"02",
          9664 => x"01",
          9665 => x"68",
          9666 => x"6f",
          9667 => x"68",
          9668 => x"00",
          9669 => x"21",
          9670 => x"25",
          9671 => x"75",
          9672 => x"73",
          9673 => x"46",
          9674 => x"65",
          9675 => x"6f",
          9676 => x"73",
          9677 => x"74",
          9678 => x"68",
          9679 => x"6f",
          9680 => x"66",
          9681 => x"20",
          9682 => x"45",
          9683 => x"00",
          9684 => x"43",
          9685 => x"6f",
          9686 => x"70",
          9687 => x"63",
          9688 => x"74",
          9689 => x"69",
          9690 => x"72",
          9691 => x"69",
          9692 => x"20",
          9693 => x"61",
          9694 => x"6e",
          9695 => x"53",
          9696 => x"22",
          9697 => x"3a",
          9698 => x"3e",
          9699 => x"7c",
          9700 => x"46",
          9701 => x"46",
          9702 => x"32",
          9703 => x"eb",
          9704 => x"53",
          9705 => x"35",
          9706 => x"4e",
          9707 => x"41",
          9708 => x"20",
          9709 => x"41",
          9710 => x"20",
          9711 => x"4e",
          9712 => x"41",
          9713 => x"20",
          9714 => x"41",
          9715 => x"20",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"80",
          9721 => x"8e",
          9722 => x"45",
          9723 => x"49",
          9724 => x"90",
          9725 => x"99",
          9726 => x"59",
          9727 => x"9c",
          9728 => x"41",
          9729 => x"a5",
          9730 => x"a8",
          9731 => x"ac",
          9732 => x"b0",
          9733 => x"b4",
          9734 => x"b8",
          9735 => x"bc",
          9736 => x"c0",
          9737 => x"c4",
          9738 => x"c8",
          9739 => x"cc",
          9740 => x"d0",
          9741 => x"d4",
          9742 => x"d8",
          9743 => x"dc",
          9744 => x"e0",
          9745 => x"e4",
          9746 => x"e8",
          9747 => x"ec",
          9748 => x"f0",
          9749 => x"f4",
          9750 => x"f8",
          9751 => x"fc",
          9752 => x"2b",
          9753 => x"3d",
          9754 => x"5c",
          9755 => x"3c",
          9756 => x"7f",
          9757 => x"00",
          9758 => x"00",
          9759 => x"01",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"01",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"01",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"01",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"01",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"01",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"01",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"01",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"01",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"01",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"01",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"01",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"01",
          9812 => x"00",
          9813 => x"00",
          9814 => x"00",
          9815 => x"01",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"01",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"01",
          9824 => x"00",
          9825 => x"00",
          9826 => x"00",
          9827 => x"01",
          9828 => x"00",
          9829 => x"00",
          9830 => x"00",
          9831 => x"01",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"01",
          9836 => x"00",
          9837 => x"00",
          9838 => x"00",
          9839 => x"01",
          9840 => x"00",
          9841 => x"00",
          9842 => x"00",
          9843 => x"01",
          9844 => x"00",
          9845 => x"00",
          9846 => x"00",
          9847 => x"01",
          9848 => x"00",
          9849 => x"00",
          9850 => x"00",
          9851 => x"01",
          9852 => x"00",
          9853 => x"00",
          9854 => x"00",
          9855 => x"01",
          9856 => x"00",
          9857 => x"00",
          9858 => x"00",
          9859 => x"01",
          9860 => x"00",
          9861 => x"00",
          9862 => x"00",
          9863 => x"01",
          9864 => x"00",
          9865 => x"00",
          9866 => x"00",
          9867 => x"01",
          9868 => x"00",
          9869 => x"00",
          9870 => x"00",
          9871 => x"00",
          9872 => x"00",
          9873 => x"00",
          9874 => x"00",
          9875 => x"00",
          9876 => x"00",
          9877 => x"00",
          9878 => x"00",
          9879 => x"01",
          9880 => x"01",
          9881 => x"00",
          9882 => x"00",
          9883 => x"00",
          9884 => x"00",
          9885 => x"05",
          9886 => x"05",
          9887 => x"05",
          9888 => x"00",
          9889 => x"01",
          9890 => x"01",
          9891 => x"01",
          9892 => x"01",
          9893 => x"00",
          9894 => x"00",
          9895 => x"00",
          9896 => x"00",
          9897 => x"00",
          9898 => x"00",
          9899 => x"00",
          9900 => x"00",
          9901 => x"00",
          9902 => x"00",
          9903 => x"00",
          9904 => x"00",
          9905 => x"00",
          9906 => x"00",
          9907 => x"00",
          9908 => x"00",
          9909 => x"00",
          9910 => x"00",
          9911 => x"00",
          9912 => x"00",
          9913 => x"00",
          9914 => x"00",
          9915 => x"00",
          9916 => x"00",
          9917 => x"00",
          9918 => x"01",
          9919 => x"00",
          9920 => x"01",
          9921 => x"00",
          9922 => x"02",
          9923 => x"00",
          9924 => x"00",
          9925 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
