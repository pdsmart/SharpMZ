zOS_BootROM.vhd