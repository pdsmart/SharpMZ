zOS_DualPortBootBRAM.vhd