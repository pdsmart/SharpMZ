-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"ff",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"92",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"e2",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"e7",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"99",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"9b",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"f8",
           386 => x"8c",
           387 => x"f8",
           388 => x"90",
           389 => x"f8",
           390 => x"8e",
           391 => x"f8",
           392 => x"90",
           393 => x"f8",
           394 => x"cd",
           395 => x"f8",
           396 => x"90",
           397 => x"f8",
           398 => x"eb",
           399 => x"f8",
           400 => x"90",
           401 => x"f8",
           402 => x"b5",
           403 => x"f8",
           404 => x"90",
           405 => x"f8",
           406 => x"b6",
           407 => x"f8",
           408 => x"90",
           409 => x"f8",
           410 => x"8e",
           411 => x"f8",
           412 => x"90",
           413 => x"f8",
           414 => x"d3",
           415 => x"f8",
           416 => x"90",
           417 => x"f8",
           418 => x"cf",
           419 => x"f8",
           420 => x"90",
           421 => x"f8",
           422 => x"db",
           423 => x"f8",
           424 => x"90",
           425 => x"f8",
           426 => x"c0",
           427 => x"f8",
           428 => x"90",
           429 => x"f8",
           430 => x"f1",
           431 => x"f8",
           432 => x"90",
           433 => x"f8",
           434 => x"95",
           435 => x"f8",
           436 => x"90",
           437 => x"f8",
           438 => x"95",
           439 => x"f8",
           440 => x"90",
           441 => x"f8",
           442 => x"e4",
           443 => x"f8",
           444 => x"90",
           445 => x"f8",
           446 => x"2d",
           447 => x"08",
           448 => x"04",
           449 => x"0c",
           450 => x"82",
           451 => x"82",
           452 => x"82",
           453 => x"be",
           454 => x"85",
           455 => x"a0",
           456 => x"85",
           457 => x"aa",
           458 => x"85",
           459 => x"a0",
           460 => x"85",
           461 => x"b7",
           462 => x"85",
           463 => x"a0",
           464 => x"85",
           465 => x"af",
           466 => x"85",
           467 => x"a0",
           468 => x"85",
           469 => x"b2",
           470 => x"85",
           471 => x"a0",
           472 => x"85",
           473 => x"bc",
           474 => x"85",
           475 => x"a0",
           476 => x"85",
           477 => x"c5",
           478 => x"85",
           479 => x"a0",
           480 => x"85",
           481 => x"b6",
           482 => x"85",
           483 => x"a0",
           484 => x"85",
           485 => x"bf",
           486 => x"85",
           487 => x"a0",
           488 => x"85",
           489 => x"c0",
           490 => x"85",
           491 => x"a0",
           492 => x"85",
           493 => x"c1",
           494 => x"85",
           495 => x"a0",
           496 => x"85",
           497 => x"c9",
           498 => x"85",
           499 => x"a0",
           500 => x"85",
           501 => x"c6",
           502 => x"85",
           503 => x"a0",
           504 => x"85",
           505 => x"cb",
           506 => x"85",
           507 => x"a0",
           508 => x"85",
           509 => x"c2",
           510 => x"85",
           511 => x"a0",
           512 => x"85",
           513 => x"ce",
           514 => x"85",
           515 => x"a0",
           516 => x"85",
           517 => x"cf",
           518 => x"85",
           519 => x"a0",
           520 => x"85",
           521 => x"b8",
           522 => x"85",
           523 => x"a0",
           524 => x"85",
           525 => x"b7",
           526 => x"85",
           527 => x"a0",
           528 => x"85",
           529 => x"b9",
           530 => x"85",
           531 => x"a0",
           532 => x"85",
           533 => x"c2",
           534 => x"85",
           535 => x"a0",
           536 => x"85",
           537 => x"d0",
           538 => x"85",
           539 => x"a0",
           540 => x"85",
           541 => x"d2",
           542 => x"85",
           543 => x"a0",
           544 => x"85",
           545 => x"d6",
           546 => x"85",
           547 => x"a0",
           548 => x"85",
           549 => x"a9",
           550 => x"85",
           551 => x"a0",
           552 => x"85",
           553 => x"d9",
           554 => x"85",
           555 => x"a0",
           556 => x"85",
           557 => x"e7",
           558 => x"85",
           559 => x"a0",
           560 => x"85",
           561 => x"e5",
           562 => x"85",
           563 => x"a0",
           564 => x"85",
           565 => x"fa",
           566 => x"85",
           567 => x"a0",
           568 => x"85",
           569 => x"fc",
           570 => x"85",
           571 => x"a0",
           572 => x"85",
           573 => x"fe",
           574 => x"85",
           575 => x"a0",
           576 => x"85",
           577 => x"ed",
           578 => x"f8",
           579 => x"90",
           580 => x"f8",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"0c",
           589 => x"82",
           590 => x"82",
           591 => x"3c",
           592 => x"10",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"10",
           598 => x"10",
           599 => x"10",
           600 => x"51",
           601 => x"73",
           602 => x"73",
           603 => x"81",
           604 => x"10",
           605 => x"07",
           606 => x"0c",
           607 => x"72",
           608 => x"81",
           609 => x"09",
           610 => x"71",
           611 => x"0a",
           612 => x"72",
           613 => x"51",
           614 => x"82",
           615 => x"82",
           616 => x"8e",
           617 => x"70",
           618 => x"0c",
           619 => x"93",
           620 => x"81",
           621 => x"04",
           622 => x"f8",
           623 => x"85",
           624 => x"3d",
           625 => x"f8",
           626 => x"08",
           627 => x"08",
           628 => x"82",
           629 => x"fc",
           630 => x"71",
           631 => x"f8",
           632 => x"08",
           633 => x"85",
           634 => x"05",
           635 => x"ff",
           636 => x"70",
           637 => x"38",
           638 => x"85",
           639 => x"05",
           640 => x"82",
           641 => x"fc",
           642 => x"85",
           643 => x"05",
           644 => x"f8",
           645 => x"08",
           646 => x"85",
           647 => x"84",
           648 => x"85",
           649 => x"82",
           650 => x"02",
           651 => x"0c",
           652 => x"82",
           653 => x"88",
           654 => x"85",
           655 => x"05",
           656 => x"f8",
           657 => x"08",
           658 => x"82",
           659 => x"8c",
           660 => x"05",
           661 => x"08",
           662 => x"82",
           663 => x"fc",
           664 => x"51",
           665 => x"82",
           666 => x"fc",
           667 => x"05",
           668 => x"08",
           669 => x"70",
           670 => x"51",
           671 => x"84",
           672 => x"39",
           673 => x"08",
           674 => x"70",
           675 => x"0c",
           676 => x"0d",
           677 => x"0c",
           678 => x"f8",
           679 => x"85",
           680 => x"3d",
           681 => x"f8",
           682 => x"08",
           683 => x"08",
           684 => x"82",
           685 => x"8c",
           686 => x"85",
           687 => x"05",
           688 => x"f8",
           689 => x"08",
           690 => x"e5",
           691 => x"f8",
           692 => x"08",
           693 => x"85",
           694 => x"05",
           695 => x"f8",
           696 => x"08",
           697 => x"85",
           698 => x"05",
           699 => x"f8",
           700 => x"08",
           701 => x"38",
           702 => x"08",
           703 => x"51",
           704 => x"85",
           705 => x"05",
           706 => x"82",
           707 => x"f8",
           708 => x"85",
           709 => x"05",
           710 => x"71",
           711 => x"85",
           712 => x"05",
           713 => x"82",
           714 => x"fc",
           715 => x"ad",
           716 => x"f8",
           717 => x"08",
           718 => x"ec",
           719 => x"3d",
           720 => x"f8",
           721 => x"85",
           722 => x"82",
           723 => x"fd",
           724 => x"85",
           725 => x"05",
           726 => x"81",
           727 => x"85",
           728 => x"05",
           729 => x"33",
           730 => x"08",
           731 => x"81",
           732 => x"f8",
           733 => x"0c",
           734 => x"08",
           735 => x"70",
           736 => x"ff",
           737 => x"54",
           738 => x"2e",
           739 => x"ce",
           740 => x"f8",
           741 => x"08",
           742 => x"82",
           743 => x"88",
           744 => x"05",
           745 => x"08",
           746 => x"70",
           747 => x"51",
           748 => x"38",
           749 => x"85",
           750 => x"05",
           751 => x"39",
           752 => x"08",
           753 => x"ff",
           754 => x"f8",
           755 => x"0c",
           756 => x"08",
           757 => x"80",
           758 => x"ff",
           759 => x"85",
           760 => x"05",
           761 => x"80",
           762 => x"85",
           763 => x"05",
           764 => x"52",
           765 => x"38",
           766 => x"85",
           767 => x"05",
           768 => x"39",
           769 => x"08",
           770 => x"ff",
           771 => x"f8",
           772 => x"0c",
           773 => x"08",
           774 => x"70",
           775 => x"70",
           776 => x"0b",
           777 => x"08",
           778 => x"ae",
           779 => x"f8",
           780 => x"08",
           781 => x"85",
           782 => x"05",
           783 => x"72",
           784 => x"82",
           785 => x"fc",
           786 => x"55",
           787 => x"8a",
           788 => x"82",
           789 => x"fc",
           790 => x"85",
           791 => x"05",
           792 => x"ec",
           793 => x"0d",
           794 => x"0c",
           795 => x"f8",
           796 => x"85",
           797 => x"3d",
           798 => x"f8",
           799 => x"08",
           800 => x"08",
           801 => x"82",
           802 => x"90",
           803 => x"2e",
           804 => x"82",
           805 => x"90",
           806 => x"05",
           807 => x"08",
           808 => x"82",
           809 => x"90",
           810 => x"05",
           811 => x"08",
           812 => x"82",
           813 => x"90",
           814 => x"2e",
           815 => x"85",
           816 => x"05",
           817 => x"82",
           818 => x"fc",
           819 => x"52",
           820 => x"82",
           821 => x"fc",
           822 => x"05",
           823 => x"08",
           824 => x"ff",
           825 => x"85",
           826 => x"05",
           827 => x"85",
           828 => x"84",
           829 => x"85",
           830 => x"82",
           831 => x"02",
           832 => x"0c",
           833 => x"80",
           834 => x"f8",
           835 => x"0c",
           836 => x"08",
           837 => x"80",
           838 => x"82",
           839 => x"88",
           840 => x"82",
           841 => x"88",
           842 => x"0b",
           843 => x"08",
           844 => x"82",
           845 => x"fc",
           846 => x"38",
           847 => x"85",
           848 => x"05",
           849 => x"f8",
           850 => x"08",
           851 => x"08",
           852 => x"82",
           853 => x"8c",
           854 => x"25",
           855 => x"85",
           856 => x"05",
           857 => x"85",
           858 => x"05",
           859 => x"82",
           860 => x"f0",
           861 => x"85",
           862 => x"05",
           863 => x"81",
           864 => x"f8",
           865 => x"0c",
           866 => x"08",
           867 => x"82",
           868 => x"fc",
           869 => x"53",
           870 => x"08",
           871 => x"52",
           872 => x"08",
           873 => x"51",
           874 => x"82",
           875 => x"70",
           876 => x"08",
           877 => x"54",
           878 => x"08",
           879 => x"80",
           880 => x"82",
           881 => x"f8",
           882 => x"82",
           883 => x"f8",
           884 => x"85",
           885 => x"05",
           886 => x"85",
           887 => x"89",
           888 => x"85",
           889 => x"82",
           890 => x"02",
           891 => x"0c",
           892 => x"80",
           893 => x"f8",
           894 => x"0c",
           895 => x"08",
           896 => x"80",
           897 => x"82",
           898 => x"88",
           899 => x"82",
           900 => x"88",
           901 => x"0b",
           902 => x"08",
           903 => x"82",
           904 => x"8c",
           905 => x"25",
           906 => x"85",
           907 => x"05",
           908 => x"85",
           909 => x"05",
           910 => x"82",
           911 => x"8c",
           912 => x"82",
           913 => x"88",
           914 => x"82",
           915 => x"85",
           916 => x"82",
           917 => x"f8",
           918 => x"82",
           919 => x"fc",
           920 => x"2e",
           921 => x"85",
           922 => x"05",
           923 => x"85",
           924 => x"05",
           925 => x"f8",
           926 => x"08",
           927 => x"ec",
           928 => x"3d",
           929 => x"f8",
           930 => x"85",
           931 => x"82",
           932 => x"ff",
           933 => x"0b",
           934 => x"08",
           935 => x"82",
           936 => x"88",
           937 => x"06",
           938 => x"09",
           939 => x"f8",
           940 => x"08",
           941 => x"f8",
           942 => x"08",
           943 => x"f8",
           944 => x"0c",
           945 => x"08",
           946 => x"81",
           947 => x"f8",
           948 => x"0c",
           949 => x"08",
           950 => x"10",
           951 => x"08",
           952 => x"51",
           953 => x"82",
           954 => x"88",
           955 => x"2e",
           956 => x"ab",
           957 => x"f8",
           958 => x"08",
           959 => x"ec",
           960 => x"3d",
           961 => x"f8",
           962 => x"85",
           963 => x"82",
           964 => x"fd",
           965 => x"53",
           966 => x"08",
           967 => x"52",
           968 => x"08",
           969 => x"51",
           970 => x"82",
           971 => x"70",
           972 => x"0c",
           973 => x"0d",
           974 => x"0c",
           975 => x"f8",
           976 => x"85",
           977 => x"3d",
           978 => x"82",
           979 => x"8c",
           980 => x"82",
           981 => x"88",
           982 => x"93",
           983 => x"ec",
           984 => x"85",
           985 => x"85",
           986 => x"85",
           987 => x"82",
           988 => x"02",
           989 => x"0c",
           990 => x"81",
           991 => x"f8",
           992 => x"0c",
           993 => x"85",
           994 => x"05",
           995 => x"f8",
           996 => x"08",
           997 => x"08",
           998 => x"27",
           999 => x"85",
          1000 => x"05",
          1001 => x"ae",
          1002 => x"82",
          1003 => x"8c",
          1004 => x"a2",
          1005 => x"f8",
          1006 => x"08",
          1007 => x"f8",
          1008 => x"0c",
          1009 => x"08",
          1010 => x"10",
          1011 => x"08",
          1012 => x"ff",
          1013 => x"85",
          1014 => x"05",
          1015 => x"80",
          1016 => x"85",
          1017 => x"05",
          1018 => x"f8",
          1019 => x"08",
          1020 => x"82",
          1021 => x"88",
          1022 => x"85",
          1023 => x"05",
          1024 => x"85",
          1025 => x"05",
          1026 => x"f8",
          1027 => x"08",
          1028 => x"08",
          1029 => x"07",
          1030 => x"08",
          1031 => x"82",
          1032 => x"fc",
          1033 => x"2a",
          1034 => x"08",
          1035 => x"82",
          1036 => x"8c",
          1037 => x"2a",
          1038 => x"08",
          1039 => x"ff",
          1040 => x"85",
          1041 => x"05",
          1042 => x"93",
          1043 => x"f8",
          1044 => x"08",
          1045 => x"f8",
          1046 => x"0c",
          1047 => x"82",
          1048 => x"f8",
          1049 => x"82",
          1050 => x"f4",
          1051 => x"82",
          1052 => x"f4",
          1053 => x"85",
          1054 => x"3d",
          1055 => x"f8",
          1056 => x"3d",
          1057 => x"08",
          1058 => x"58",
          1059 => x"80",
          1060 => x"39",
          1061 => x"f2",
          1062 => x"85",
          1063 => x"78",
          1064 => x"33",
          1065 => x"39",
          1066 => x"73",
          1067 => x"81",
          1068 => x"81",
          1069 => x"39",
          1070 => x"84",
          1071 => x"ec",
          1072 => x"52",
          1073 => x"3f",
          1074 => x"08",
          1075 => x"75",
          1076 => x"f2",
          1077 => x"ec",
          1078 => x"84",
          1079 => x"73",
          1080 => x"b0",
          1081 => x"70",
          1082 => x"58",
          1083 => x"27",
          1084 => x"54",
          1085 => x"ec",
          1086 => x"0d",
          1087 => x"0d",
          1088 => x"93",
          1089 => x"38",
          1090 => x"52",
          1091 => x"12",
          1092 => x"ea",
          1093 => x"80",
          1094 => x"80",
          1095 => x"39",
          1096 => x"51",
          1097 => x"81",
          1098 => x"80",
          1099 => x"eb",
          1100 => x"e4",
          1101 => x"c8",
          1102 => x"39",
          1103 => x"51",
          1104 => x"81",
          1105 => x"80",
          1106 => x"ec",
          1107 => x"c8",
          1108 => x"9c",
          1109 => x"39",
          1110 => x"51",
          1111 => x"ec",
          1112 => x"39",
          1113 => x"51",
          1114 => x"ed",
          1115 => x"39",
          1116 => x"51",
          1117 => x"ed",
          1118 => x"39",
          1119 => x"51",
          1120 => x"ed",
          1121 => x"39",
          1122 => x"51",
          1123 => x"ee",
          1124 => x"39",
          1125 => x"51",
          1126 => x"83",
          1127 => x"fb",
          1128 => x"79",
          1129 => x"87",
          1130 => x"38",
          1131 => x"75",
          1132 => x"3f",
          1133 => x"85",
          1134 => x"90",
          1135 => x"52",
          1136 => x"c6",
          1137 => x"ec",
          1138 => x"51",
          1139 => x"82",
          1140 => x"54",
          1141 => x"52",
          1142 => x"51",
          1143 => x"87",
          1144 => x"ec",
          1145 => x"02",
          1146 => x"e3",
          1147 => x"57",
          1148 => x"09",
          1149 => x"7a",
          1150 => x"51",
          1151 => x"78",
          1152 => x"ff",
          1153 => x"81",
          1154 => x"07",
          1155 => x"06",
          1156 => x"56",
          1157 => x"38",
          1158 => x"52",
          1159 => x"52",
          1160 => x"98",
          1161 => x"ec",
          1162 => x"85",
          1163 => x"38",
          1164 => x"08",
          1165 => x"88",
          1166 => x"ec",
          1167 => x"3d",
          1168 => x"84",
          1169 => x"52",
          1170 => x"8a",
          1171 => x"85",
          1172 => x"82",
          1173 => x"90",
          1174 => x"74",
          1175 => x"38",
          1176 => x"19",
          1177 => x"39",
          1178 => x"05",
          1179 => x"bf",
          1180 => x"81",
          1181 => x"07",
          1182 => x"09",
          1183 => x"9f",
          1184 => x"51",
          1185 => x"74",
          1186 => x"38",
          1187 => x"53",
          1188 => x"88",
          1189 => x"51",
          1190 => x"76",
          1191 => x"85",
          1192 => x"3d",
          1193 => x"3d",
          1194 => x"84",
          1195 => x"33",
          1196 => x"57",
          1197 => x"52",
          1198 => x"a7",
          1199 => x"ec",
          1200 => x"75",
          1201 => x"38",
          1202 => x"98",
          1203 => x"60",
          1204 => x"82",
          1205 => x"7e",
          1206 => x"77",
          1207 => x"ec",
          1208 => x"39",
          1209 => x"82",
          1210 => x"89",
          1211 => x"f3",
          1212 => x"61",
          1213 => x"05",
          1214 => x"33",
          1215 => x"68",
          1216 => x"5c",
          1217 => x"7a",
          1218 => x"e8",
          1219 => x"3f",
          1220 => x"51",
          1221 => x"80",
          1222 => x"27",
          1223 => x"7b",
          1224 => x"38",
          1225 => x"a4",
          1226 => x"39",
          1227 => x"72",
          1228 => x"38",
          1229 => x"81",
          1230 => x"ae",
          1231 => x"39",
          1232 => x"51",
          1233 => x"82",
          1234 => x"39",
          1235 => x"72",
          1236 => x"38",
          1237 => x"81",
          1238 => x"ad",
          1239 => x"39",
          1240 => x"51",
          1241 => x"84",
          1242 => x"39",
          1243 => x"72",
          1244 => x"38",
          1245 => x"81",
          1246 => x"ad",
          1247 => x"39",
          1248 => x"51",
          1249 => x"81",
          1250 => x"51",
          1251 => x"ff",
          1252 => x"ef",
          1253 => x"d3",
          1254 => x"74",
          1255 => x"38",
          1256 => x"33",
          1257 => x"56",
          1258 => x"83",
          1259 => x"80",
          1260 => x"27",
          1261 => x"53",
          1262 => x"70",
          1263 => x"51",
          1264 => x"2e",
          1265 => x"80",
          1266 => x"38",
          1267 => x"39",
          1268 => x"ba",
          1269 => x"55",
          1270 => x"ef",
          1271 => x"8b",
          1272 => x"79",
          1273 => x"9b",
          1274 => x"85",
          1275 => x"2b",
          1276 => x"51",
          1277 => x"2e",
          1278 => x"ae",
          1279 => x"3f",
          1280 => x"08",
          1281 => x"98",
          1282 => x"32",
          1283 => x"05",
          1284 => x"70",
          1285 => x"70",
          1286 => x"75",
          1287 => x"58",
          1288 => x"51",
          1289 => x"24",
          1290 => x"9b",
          1291 => x"06",
          1292 => x"53",
          1293 => x"1e",
          1294 => x"26",
          1295 => x"ff",
          1296 => x"85",
          1297 => x"3d",
          1298 => x"3d",
          1299 => x"05",
          1300 => x"9c",
          1301 => x"a0",
          1302 => x"ff",
          1303 => x"c4",
          1304 => x"d1",
          1305 => x"ac",
          1306 => x"b8",
          1307 => x"c5",
          1308 => x"ef",
          1309 => x"e3",
          1310 => x"2e",
          1311 => x"86",
          1312 => x"0d",
          1313 => x"0d",
          1314 => x"80",
          1315 => x"ec",
          1316 => x"96",
          1317 => x"ef",
          1318 => x"e0",
          1319 => x"96",
          1320 => x"81",
          1321 => x"06",
          1322 => x"80",
          1323 => x"81",
          1324 => x"3f",
          1325 => x"51",
          1326 => x"80",
          1327 => x"3f",
          1328 => x"70",
          1329 => x"52",
          1330 => x"92",
          1331 => x"96",
          1332 => x"f0",
          1333 => x"a4",
          1334 => x"96",
          1335 => x"83",
          1336 => x"06",
          1337 => x"80",
          1338 => x"81",
          1339 => x"3f",
          1340 => x"51",
          1341 => x"80",
          1342 => x"3f",
          1343 => x"70",
          1344 => x"52",
          1345 => x"92",
          1346 => x"95",
          1347 => x"f0",
          1348 => x"e8",
          1349 => x"95",
          1350 => x"85",
          1351 => x"06",
          1352 => x"80",
          1353 => x"81",
          1354 => x"3f",
          1355 => x"51",
          1356 => x"80",
          1357 => x"3f",
          1358 => x"70",
          1359 => x"52",
          1360 => x"92",
          1361 => x"95",
          1362 => x"f0",
          1363 => x"ac",
          1364 => x"95",
          1365 => x"87",
          1366 => x"06",
          1367 => x"80",
          1368 => x"81",
          1369 => x"3f",
          1370 => x"51",
          1371 => x"80",
          1372 => x"3f",
          1373 => x"70",
          1374 => x"52",
          1375 => x"92",
          1376 => x"94",
          1377 => x"f0",
          1378 => x"f0",
          1379 => x"94",
          1380 => x"f0",
          1381 => x"0d",
          1382 => x"0d",
          1383 => x"05",
          1384 => x"70",
          1385 => x"80",
          1386 => x"ed",
          1387 => x"0b",
          1388 => x"33",
          1389 => x"38",
          1390 => x"f1",
          1391 => x"9c",
          1392 => x"fe",
          1393 => x"85",
          1394 => x"81",
          1395 => x"85",
          1396 => x"80",
          1397 => x"31",
          1398 => x"73",
          1399 => x"80",
          1400 => x"0b",
          1401 => x"33",
          1402 => x"2e",
          1403 => x"af",
          1404 => x"cc",
          1405 => x"75",
          1406 => x"c4",
          1407 => x"ec",
          1408 => x"8b",
          1409 => x"ec",
          1410 => x"df",
          1411 => x"82",
          1412 => x"81",
          1413 => x"82",
          1414 => x"82",
          1415 => x"0b",
          1416 => x"e8",
          1417 => x"82",
          1418 => x"06",
          1419 => x"f1",
          1420 => x"52",
          1421 => x"92",
          1422 => x"82",
          1423 => x"87",
          1424 => x"ce",
          1425 => x"70",
          1426 => x"c8",
          1427 => x"81",
          1428 => x"80",
          1429 => x"82",
          1430 => x"81",
          1431 => x"78",
          1432 => x"81",
          1433 => x"81",
          1434 => x"96",
          1435 => x"59",
          1436 => x"7c",
          1437 => x"82",
          1438 => x"80",
          1439 => x"82",
          1440 => x"7d",
          1441 => x"81",
          1442 => x"8d",
          1443 => x"70",
          1444 => x"f2",
          1445 => x"d3",
          1446 => x"70",
          1447 => x"f8",
          1448 => x"fd",
          1449 => x"3d",
          1450 => x"51",
          1451 => x"82",
          1452 => x"90",
          1453 => x"2c",
          1454 => x"80",
          1455 => x"9c",
          1456 => x"c2",
          1457 => x"78",
          1458 => x"d1",
          1459 => x"24",
          1460 => x"80",
          1461 => x"38",
          1462 => x"80",
          1463 => x"bb",
          1464 => x"c0",
          1465 => x"38",
          1466 => x"24",
          1467 => x"78",
          1468 => x"8a",
          1469 => x"39",
          1470 => x"2e",
          1471 => x"78",
          1472 => x"92",
          1473 => x"c3",
          1474 => x"38",
          1475 => x"2e",
          1476 => x"8a",
          1477 => x"81",
          1478 => x"ed",
          1479 => x"83",
          1480 => x"78",
          1481 => x"89",
          1482 => x"ef",
          1483 => x"85",
          1484 => x"38",
          1485 => x"b4",
          1486 => x"11",
          1487 => x"05",
          1488 => x"3f",
          1489 => x"08",
          1490 => x"c6",
          1491 => x"fe",
          1492 => x"ff",
          1493 => x"a7",
          1494 => x"85",
          1495 => x"2e",
          1496 => x"b4",
          1497 => x"11",
          1498 => x"05",
          1499 => x"3f",
          1500 => x"08",
          1501 => x"85",
          1502 => x"81",
          1503 => x"9f",
          1504 => x"63",
          1505 => x"7b",
          1506 => x"38",
          1507 => x"7a",
          1508 => x"5c",
          1509 => x"26",
          1510 => x"d8",
          1511 => x"ff",
          1512 => x"ff",
          1513 => x"a7",
          1514 => x"85",
          1515 => x"2e",
          1516 => x"b4",
          1517 => x"11",
          1518 => x"05",
          1519 => x"3f",
          1520 => x"08",
          1521 => x"ca",
          1522 => x"fe",
          1523 => x"ff",
          1524 => x"a6",
          1525 => x"85",
          1526 => x"2e",
          1527 => x"81",
          1528 => x"9f",
          1529 => x"5a",
          1530 => x"81",
          1531 => x"59",
          1532 => x"05",
          1533 => x"34",
          1534 => x"42",
          1535 => x"3d",
          1536 => x"53",
          1537 => x"51",
          1538 => x"82",
          1539 => x"80",
          1540 => x"38",
          1541 => x"fc",
          1542 => x"84",
          1543 => x"b3",
          1544 => x"ec",
          1545 => x"fc",
          1546 => x"3d",
          1547 => x"53",
          1548 => x"51",
          1549 => x"82",
          1550 => x"80",
          1551 => x"38",
          1552 => x"51",
          1553 => x"63",
          1554 => x"27",
          1555 => x"70",
          1556 => x"5e",
          1557 => x"7c",
          1558 => x"78",
          1559 => x"79",
          1560 => x"52",
          1561 => x"51",
          1562 => x"81",
          1563 => x"05",
          1564 => x"39",
          1565 => x"51",
          1566 => x"b4",
          1567 => x"11",
          1568 => x"05",
          1569 => x"3f",
          1570 => x"08",
          1571 => x"82",
          1572 => x"59",
          1573 => x"89",
          1574 => x"90",
          1575 => x"cd",
          1576 => x"d9",
          1577 => x"80",
          1578 => x"82",
          1579 => x"44",
          1580 => x"84",
          1581 => x"78",
          1582 => x"38",
          1583 => x"08",
          1584 => x"82",
          1585 => x"59",
          1586 => x"88",
          1587 => x"a8",
          1588 => x"39",
          1589 => x"33",
          1590 => x"2e",
          1591 => x"84",
          1592 => x"89",
          1593 => x"c0",
          1594 => x"05",
          1595 => x"fe",
          1596 => x"ff",
          1597 => x"a4",
          1598 => x"85",
          1599 => x"de",
          1600 => x"d8",
          1601 => x"80",
          1602 => x"82",
          1603 => x"43",
          1604 => x"82",
          1605 => x"59",
          1606 => x"88",
          1607 => x"9c",
          1608 => x"39",
          1609 => x"33",
          1610 => x"2e",
          1611 => x"84",
          1612 => x"aa",
          1613 => x"db",
          1614 => x"80",
          1615 => x"82",
          1616 => x"43",
          1617 => x"84",
          1618 => x"78",
          1619 => x"38",
          1620 => x"08",
          1621 => x"82",
          1622 => x"88",
          1623 => x"3d",
          1624 => x"53",
          1625 => x"51",
          1626 => x"82",
          1627 => x"80",
          1628 => x"80",
          1629 => x"7a",
          1630 => x"38",
          1631 => x"90",
          1632 => x"81",
          1633 => x"07",
          1634 => x"7f",
          1635 => x"5a",
          1636 => x"2e",
          1637 => x"a0",
          1638 => x"88",
          1639 => x"dc",
          1640 => x"3f",
          1641 => x"54",
          1642 => x"52",
          1643 => x"bf",
          1644 => x"ec",
          1645 => x"3f",
          1646 => x"b4",
          1647 => x"11",
          1648 => x"05",
          1649 => x"3f",
          1650 => x"08",
          1651 => x"c2",
          1652 => x"fe",
          1653 => x"ff",
          1654 => x"a2",
          1655 => x"85",
          1656 => x"2e",
          1657 => x"59",
          1658 => x"05",
          1659 => x"63",
          1660 => x"b4",
          1661 => x"11",
          1662 => x"05",
          1663 => x"3f",
          1664 => x"08",
          1665 => x"8a",
          1666 => x"33",
          1667 => x"f2",
          1668 => x"c7",
          1669 => x"52",
          1670 => x"99",
          1671 => x"79",
          1672 => x"ae",
          1673 => x"38",
          1674 => x"9f",
          1675 => x"fe",
          1676 => x"ff",
          1677 => x"a2",
          1678 => x"85",
          1679 => x"2e",
          1680 => x"59",
          1681 => x"05",
          1682 => x"63",
          1683 => x"ff",
          1684 => x"f3",
          1685 => x"93",
          1686 => x"39",
          1687 => x"f4",
          1688 => x"84",
          1689 => x"e7",
          1690 => x"ec",
          1691 => x"f8",
          1692 => x"3d",
          1693 => x"53",
          1694 => x"51",
          1695 => x"82",
          1696 => x"80",
          1697 => x"60",
          1698 => x"05",
          1699 => x"82",
          1700 => x"78",
          1701 => x"fe",
          1702 => x"ff",
          1703 => x"a3",
          1704 => x"85",
          1705 => x"38",
          1706 => x"60",
          1707 => x"52",
          1708 => x"51",
          1709 => x"80",
          1710 => x"51",
          1711 => x"79",
          1712 => x"59",
          1713 => x"f7",
          1714 => x"9f",
          1715 => x"60",
          1716 => x"d7",
          1717 => x"fe",
          1718 => x"ff",
          1719 => x"a2",
          1720 => x"85",
          1721 => x"2e",
          1722 => x"59",
          1723 => x"22",
          1724 => x"05",
          1725 => x"41",
          1726 => x"81",
          1727 => x"98",
          1728 => x"a7",
          1729 => x"fe",
          1730 => x"ff",
          1731 => x"a2",
          1732 => x"85",
          1733 => x"2e",
          1734 => x"b4",
          1735 => x"11",
          1736 => x"05",
          1737 => x"3f",
          1738 => x"08",
          1739 => x"38",
          1740 => x"0c",
          1741 => x"05",
          1742 => x"fe",
          1743 => x"ff",
          1744 => x"a2",
          1745 => x"85",
          1746 => x"38",
          1747 => x"60",
          1748 => x"52",
          1749 => x"51",
          1750 => x"80",
          1751 => x"51",
          1752 => x"79",
          1753 => x"59",
          1754 => x"f6",
          1755 => x"79",
          1756 => x"b4",
          1757 => x"11",
          1758 => x"05",
          1759 => x"3f",
          1760 => x"08",
          1761 => x"38",
          1762 => x"0c",
          1763 => x"05",
          1764 => x"39",
          1765 => x"51",
          1766 => x"ff",
          1767 => x"3d",
          1768 => x"53",
          1769 => x"51",
          1770 => x"82",
          1771 => x"80",
          1772 => x"38",
          1773 => x"f3",
          1774 => x"9f",
          1775 => x"78",
          1776 => x"ff",
          1777 => x"ff",
          1778 => x"9f",
          1779 => x"85",
          1780 => x"2e",
          1781 => x"63",
          1782 => x"c0",
          1783 => x"3f",
          1784 => x"2d",
          1785 => x"08",
          1786 => x"a6",
          1787 => x"ec",
          1788 => x"f3",
          1789 => x"e3",
          1790 => x"39",
          1791 => x"51",
          1792 => x"db",
          1793 => x"8a",
          1794 => x"94",
          1795 => x"3f",
          1796 => x"ab",
          1797 => x"3f",
          1798 => x"79",
          1799 => x"59",
          1800 => x"f4",
          1801 => x"7d",
          1802 => x"80",
          1803 => x"38",
          1804 => x"84",
          1805 => x"b5",
          1806 => x"ec",
          1807 => x"5b",
          1808 => x"b1",
          1809 => x"24",
          1810 => x"81",
          1811 => x"80",
          1812 => x"83",
          1813 => x"80",
          1814 => x"f4",
          1815 => x"55",
          1816 => x"54",
          1817 => x"f4",
          1818 => x"3d",
          1819 => x"51",
          1820 => x"b8",
          1821 => x"d0",
          1822 => x"ff",
          1823 => x"9b",
          1824 => x"39",
          1825 => x"f4",
          1826 => x"53",
          1827 => x"52",
          1828 => x"b0",
          1829 => x"d9",
          1830 => x"7b",
          1831 => x"81",
          1832 => x"b4",
          1833 => x"05",
          1834 => x"3f",
          1835 => x"58",
          1836 => x"57",
          1837 => x"55",
          1838 => x"a0",
          1839 => x"a0",
          1840 => x"3d",
          1841 => x"51",
          1842 => x"82",
          1843 => x"82",
          1844 => x"09",
          1845 => x"05",
          1846 => x"80",
          1847 => x"5b",
          1848 => x"7a",
          1849 => x"38",
          1850 => x"7a",
          1851 => x"80",
          1852 => x"81",
          1853 => x"ff",
          1854 => x"7a",
          1855 => x"7d",
          1856 => x"81",
          1857 => x"78",
          1858 => x"ff",
          1859 => x"06",
          1860 => x"81",
          1861 => x"9a",
          1862 => x"f6",
          1863 => x"0d",
          1864 => x"85",
          1865 => x"c0",
          1866 => x"08",
          1867 => x"84",
          1868 => x"51",
          1869 => x"82",
          1870 => x"90",
          1871 => x"55",
          1872 => x"80",
          1873 => x"e3",
          1874 => x"82",
          1875 => x"07",
          1876 => x"c0",
          1877 => x"08",
          1878 => x"84",
          1879 => x"51",
          1880 => x"82",
          1881 => x"90",
          1882 => x"55",
          1883 => x"80",
          1884 => x"e3",
          1885 => x"82",
          1886 => x"07",
          1887 => x"80",
          1888 => x"c0",
          1889 => x"8c",
          1890 => x"87",
          1891 => x"0c",
          1892 => x"0b",
          1893 => x"0c",
          1894 => x"0b",
          1895 => x"0c",
          1896 => x"92",
          1897 => x"f4",
          1898 => x"bf",
          1899 => x"f0",
          1900 => x"3f",
          1901 => x"92",
          1902 => x"51",
          1903 => x"f1",
          1904 => x"04",
          1905 => x"80",
          1906 => x"71",
          1907 => x"87",
          1908 => x"85",
          1909 => x"ff",
          1910 => x"ff",
          1911 => x"72",
          1912 => x"38",
          1913 => x"ec",
          1914 => x"0d",
          1915 => x"0d",
          1916 => x"54",
          1917 => x"52",
          1918 => x"2e",
          1919 => x"72",
          1920 => x"a0",
          1921 => x"06",
          1922 => x"13",
          1923 => x"72",
          1924 => x"a2",
          1925 => x"06",
          1926 => x"13",
          1927 => x"72",
          1928 => x"2e",
          1929 => x"9f",
          1930 => x"81",
          1931 => x"72",
          1932 => x"70",
          1933 => x"38",
          1934 => x"80",
          1935 => x"73",
          1936 => x"39",
          1937 => x"80",
          1938 => x"54",
          1939 => x"83",
          1940 => x"70",
          1941 => x"38",
          1942 => x"80",
          1943 => x"54",
          1944 => x"09",
          1945 => x"38",
          1946 => x"a2",
          1947 => x"81",
          1948 => x"25",
          1949 => x"51",
          1950 => x"2e",
          1951 => x"72",
          1952 => x"54",
          1953 => x"0c",
          1954 => x"82",
          1955 => x"86",
          1956 => x"fc",
          1957 => x"53",
          1958 => x"2e",
          1959 => x"3d",
          1960 => x"72",
          1961 => x"3f",
          1962 => x"08",
          1963 => x"53",
          1964 => x"53",
          1965 => x"ec",
          1966 => x"0d",
          1967 => x"0d",
          1968 => x"33",
          1969 => x"53",
          1970 => x"8b",
          1971 => x"38",
          1972 => x"ff",
          1973 => x"52",
          1974 => x"81",
          1975 => x"13",
          1976 => x"52",
          1977 => x"80",
          1978 => x"13",
          1979 => x"52",
          1980 => x"80",
          1981 => x"13",
          1982 => x"52",
          1983 => x"80",
          1984 => x"13",
          1985 => x"52",
          1986 => x"26",
          1987 => x"8a",
          1988 => x"87",
          1989 => x"e7",
          1990 => x"38",
          1991 => x"c0",
          1992 => x"72",
          1993 => x"98",
          1994 => x"13",
          1995 => x"98",
          1996 => x"13",
          1997 => x"98",
          1998 => x"13",
          1999 => x"98",
          2000 => x"13",
          2001 => x"98",
          2002 => x"13",
          2003 => x"98",
          2004 => x"87",
          2005 => x"0c",
          2006 => x"98",
          2007 => x"0b",
          2008 => x"9c",
          2009 => x"71",
          2010 => x"0c",
          2011 => x"04",
          2012 => x"7f",
          2013 => x"98",
          2014 => x"7d",
          2015 => x"98",
          2016 => x"7d",
          2017 => x"c0",
          2018 => x"5a",
          2019 => x"34",
          2020 => x"b4",
          2021 => x"83",
          2022 => x"c0",
          2023 => x"5a",
          2024 => x"34",
          2025 => x"ac",
          2026 => x"85",
          2027 => x"c0",
          2028 => x"5a",
          2029 => x"34",
          2030 => x"a4",
          2031 => x"88",
          2032 => x"c0",
          2033 => x"5a",
          2034 => x"23",
          2035 => x"79",
          2036 => x"06",
          2037 => x"ff",
          2038 => x"86",
          2039 => x"85",
          2040 => x"84",
          2041 => x"83",
          2042 => x"82",
          2043 => x"7d",
          2044 => x"06",
          2045 => x"88",
          2046 => x"3f",
          2047 => x"04",
          2048 => x"02",
          2049 => x"70",
          2050 => x"70",
          2051 => x"52",
          2052 => x"84",
          2053 => x"3d",
          2054 => x"3d",
          2055 => x"84",
          2056 => x"81",
          2057 => x"55",
          2058 => x"94",
          2059 => x"80",
          2060 => x"87",
          2061 => x"51",
          2062 => x"96",
          2063 => x"06",
          2064 => x"70",
          2065 => x"38",
          2066 => x"70",
          2067 => x"51",
          2068 => x"72",
          2069 => x"81",
          2070 => x"70",
          2071 => x"38",
          2072 => x"70",
          2073 => x"51",
          2074 => x"38",
          2075 => x"06",
          2076 => x"94",
          2077 => x"80",
          2078 => x"87",
          2079 => x"52",
          2080 => x"75",
          2081 => x"0c",
          2082 => x"04",
          2083 => x"02",
          2084 => x"82",
          2085 => x"70",
          2086 => x"57",
          2087 => x"c0",
          2088 => x"74",
          2089 => x"38",
          2090 => x"94",
          2091 => x"70",
          2092 => x"81",
          2093 => x"52",
          2094 => x"8c",
          2095 => x"2a",
          2096 => x"51",
          2097 => x"38",
          2098 => x"70",
          2099 => x"51",
          2100 => x"8d",
          2101 => x"2a",
          2102 => x"51",
          2103 => x"be",
          2104 => x"ff",
          2105 => x"c0",
          2106 => x"70",
          2107 => x"38",
          2108 => x"90",
          2109 => x"0c",
          2110 => x"04",
          2111 => x"79",
          2112 => x"33",
          2113 => x"06",
          2114 => x"70",
          2115 => x"fc",
          2116 => x"ff",
          2117 => x"82",
          2118 => x"70",
          2119 => x"59",
          2120 => x"87",
          2121 => x"51",
          2122 => x"86",
          2123 => x"94",
          2124 => x"08",
          2125 => x"70",
          2126 => x"54",
          2127 => x"2e",
          2128 => x"91",
          2129 => x"06",
          2130 => x"d7",
          2131 => x"32",
          2132 => x"51",
          2133 => x"2e",
          2134 => x"93",
          2135 => x"06",
          2136 => x"ff",
          2137 => x"81",
          2138 => x"87",
          2139 => x"52",
          2140 => x"86",
          2141 => x"94",
          2142 => x"72",
          2143 => x"74",
          2144 => x"ff",
          2145 => x"57",
          2146 => x"38",
          2147 => x"ec",
          2148 => x"0d",
          2149 => x"0d",
          2150 => x"33",
          2151 => x"06",
          2152 => x"c0",
          2153 => x"72",
          2154 => x"38",
          2155 => x"94",
          2156 => x"70",
          2157 => x"81",
          2158 => x"51",
          2159 => x"e2",
          2160 => x"ff",
          2161 => x"c0",
          2162 => x"70",
          2163 => x"38",
          2164 => x"90",
          2165 => x"70",
          2166 => x"82",
          2167 => x"51",
          2168 => x"04",
          2169 => x"82",
          2170 => x"70",
          2171 => x"52",
          2172 => x"94",
          2173 => x"80",
          2174 => x"87",
          2175 => x"52",
          2176 => x"82",
          2177 => x"06",
          2178 => x"ff",
          2179 => x"2e",
          2180 => x"81",
          2181 => x"87",
          2182 => x"52",
          2183 => x"86",
          2184 => x"94",
          2185 => x"08",
          2186 => x"70",
          2187 => x"53",
          2188 => x"85",
          2189 => x"3d",
          2190 => x"3d",
          2191 => x"9e",
          2192 => x"9c",
          2193 => x"51",
          2194 => x"2e",
          2195 => x"87",
          2196 => x"08",
          2197 => x"0c",
          2198 => x"a8",
          2199 => x"94",
          2200 => x"9e",
          2201 => x"84",
          2202 => x"c0",
          2203 => x"82",
          2204 => x"87",
          2205 => x"08",
          2206 => x"0c",
          2207 => x"a0",
          2208 => x"a4",
          2209 => x"9e",
          2210 => x"84",
          2211 => x"c0",
          2212 => x"82",
          2213 => x"87",
          2214 => x"08",
          2215 => x"0c",
          2216 => x"b8",
          2217 => x"b4",
          2218 => x"9e",
          2219 => x"84",
          2220 => x"c0",
          2221 => x"82",
          2222 => x"87",
          2223 => x"08",
          2224 => x"0c",
          2225 => x"80",
          2226 => x"82",
          2227 => x"87",
          2228 => x"08",
          2229 => x"0c",
          2230 => x"88",
          2231 => x"cc",
          2232 => x"9e",
          2233 => x"84",
          2234 => x"0b",
          2235 => x"34",
          2236 => x"c0",
          2237 => x"70",
          2238 => x"06",
          2239 => x"70",
          2240 => x"38",
          2241 => x"82",
          2242 => x"80",
          2243 => x"9e",
          2244 => x"88",
          2245 => x"51",
          2246 => x"80",
          2247 => x"81",
          2248 => x"84",
          2249 => x"0b",
          2250 => x"90",
          2251 => x"80",
          2252 => x"52",
          2253 => x"2e",
          2254 => x"52",
          2255 => x"d7",
          2256 => x"87",
          2257 => x"08",
          2258 => x"80",
          2259 => x"52",
          2260 => x"83",
          2261 => x"71",
          2262 => x"34",
          2263 => x"c0",
          2264 => x"70",
          2265 => x"06",
          2266 => x"70",
          2267 => x"38",
          2268 => x"82",
          2269 => x"80",
          2270 => x"9e",
          2271 => x"90",
          2272 => x"51",
          2273 => x"80",
          2274 => x"81",
          2275 => x"84",
          2276 => x"0b",
          2277 => x"90",
          2278 => x"80",
          2279 => x"52",
          2280 => x"2e",
          2281 => x"52",
          2282 => x"db",
          2283 => x"87",
          2284 => x"08",
          2285 => x"80",
          2286 => x"52",
          2287 => x"83",
          2288 => x"71",
          2289 => x"34",
          2290 => x"c0",
          2291 => x"70",
          2292 => x"06",
          2293 => x"70",
          2294 => x"38",
          2295 => x"82",
          2296 => x"80",
          2297 => x"9e",
          2298 => x"80",
          2299 => x"51",
          2300 => x"80",
          2301 => x"81",
          2302 => x"84",
          2303 => x"0b",
          2304 => x"90",
          2305 => x"80",
          2306 => x"52",
          2307 => x"83",
          2308 => x"71",
          2309 => x"34",
          2310 => x"90",
          2311 => x"80",
          2312 => x"2a",
          2313 => x"70",
          2314 => x"34",
          2315 => x"c0",
          2316 => x"70",
          2317 => x"51",
          2318 => x"80",
          2319 => x"81",
          2320 => x"84",
          2321 => x"c0",
          2322 => x"70",
          2323 => x"70",
          2324 => x"51",
          2325 => x"84",
          2326 => x"0b",
          2327 => x"90",
          2328 => x"06",
          2329 => x"70",
          2330 => x"38",
          2331 => x"82",
          2332 => x"87",
          2333 => x"08",
          2334 => x"51",
          2335 => x"84",
          2336 => x"3d",
          2337 => x"3d",
          2338 => x"a0",
          2339 => x"3f",
          2340 => x"33",
          2341 => x"2e",
          2342 => x"f5",
          2343 => x"cb",
          2344 => x"c8",
          2345 => x"3f",
          2346 => x"33",
          2347 => x"2e",
          2348 => x"84",
          2349 => x"84",
          2350 => x"54",
          2351 => x"e0",
          2352 => x"3f",
          2353 => x"33",
          2354 => x"2e",
          2355 => x"84",
          2356 => x"84",
          2357 => x"54",
          2358 => x"fc",
          2359 => x"3f",
          2360 => x"33",
          2361 => x"2e",
          2362 => x"84",
          2363 => x"84",
          2364 => x"54",
          2365 => x"98",
          2366 => x"3f",
          2367 => x"33",
          2368 => x"2e",
          2369 => x"84",
          2370 => x"84",
          2371 => x"54",
          2372 => x"b4",
          2373 => x"3f",
          2374 => x"33",
          2375 => x"2e",
          2376 => x"84",
          2377 => x"84",
          2378 => x"54",
          2379 => x"d0",
          2380 => x"3f",
          2381 => x"33",
          2382 => x"2e",
          2383 => x"84",
          2384 => x"81",
          2385 => x"8a",
          2386 => x"84",
          2387 => x"73",
          2388 => x"38",
          2389 => x"33",
          2390 => x"8c",
          2391 => x"3f",
          2392 => x"33",
          2393 => x"2e",
          2394 => x"84",
          2395 => x"81",
          2396 => x"89",
          2397 => x"84",
          2398 => x"73",
          2399 => x"38",
          2400 => x"51",
          2401 => x"82",
          2402 => x"54",
          2403 => x"88",
          2404 => x"e0",
          2405 => x"3f",
          2406 => x"33",
          2407 => x"2e",
          2408 => x"f7",
          2409 => x"c3",
          2410 => x"dd",
          2411 => x"80",
          2412 => x"81",
          2413 => x"83",
          2414 => x"84",
          2415 => x"73",
          2416 => x"38",
          2417 => x"51",
          2418 => x"81",
          2419 => x"83",
          2420 => x"84",
          2421 => x"81",
          2422 => x"88",
          2423 => x"84",
          2424 => x"81",
          2425 => x"88",
          2426 => x"84",
          2427 => x"81",
          2428 => x"88",
          2429 => x"f9",
          2430 => x"ef",
          2431 => x"c4",
          2432 => x"f9",
          2433 => x"d3",
          2434 => x"c8",
          2435 => x"84",
          2436 => x"51",
          2437 => x"82",
          2438 => x"54",
          2439 => x"52",
          2440 => x"08",
          2441 => x"3f",
          2442 => x"ec",
          2443 => x"73",
          2444 => x"c4",
          2445 => x"3f",
          2446 => x"33",
          2447 => x"2e",
          2448 => x"84",
          2449 => x"bd",
          2450 => x"74",
          2451 => x"3f",
          2452 => x"08",
          2453 => x"c0",
          2454 => x"ec",
          2455 => x"aa",
          2456 => x"85",
          2457 => x"53",
          2458 => x"f9",
          2459 => x"eb",
          2460 => x"d6",
          2461 => x"80",
          2462 => x"82",
          2463 => x"55",
          2464 => x"52",
          2465 => x"82",
          2466 => x"ec",
          2467 => x"84",
          2468 => x"85",
          2469 => x"cf",
          2470 => x"82",
          2471 => x"31",
          2472 => x"81",
          2473 => x"87",
          2474 => x"f2",
          2475 => x"bb",
          2476 => x"0d",
          2477 => x"0d",
          2478 => x"33",
          2479 => x"71",
          2480 => x"38",
          2481 => x"52",
          2482 => x"12",
          2483 => x"fa",
          2484 => x"39",
          2485 => x"51",
          2486 => x"fa",
          2487 => x"39",
          2488 => x"51",
          2489 => x"fa",
          2490 => x"39",
          2491 => x"51",
          2492 => x"84",
          2493 => x"71",
          2494 => x"04",
          2495 => x"c0",
          2496 => x"04",
          2497 => x"08",
          2498 => x"84",
          2499 => x"3d",
          2500 => x"05",
          2501 => x"8a",
          2502 => x"06",
          2503 => x"51",
          2504 => x"9c",
          2505 => x"71",
          2506 => x"38",
          2507 => x"82",
          2508 => x"81",
          2509 => x"fc",
          2510 => x"82",
          2511 => x"52",
          2512 => x"85",
          2513 => x"71",
          2514 => x"0d",
          2515 => x"0d",
          2516 => x"33",
          2517 => x"08",
          2518 => x"f4",
          2519 => x"ff",
          2520 => x"82",
          2521 => x"84",
          2522 => x"fd",
          2523 => x"54",
          2524 => x"81",
          2525 => x"53",
          2526 => x"8e",
          2527 => x"ff",
          2528 => x"14",
          2529 => x"3f",
          2530 => x"3d",
          2531 => x"3d",
          2532 => x"9c",
          2533 => x"82",
          2534 => x"56",
          2535 => x"70",
          2536 => x"53",
          2537 => x"2e",
          2538 => x"81",
          2539 => x"81",
          2540 => x"da",
          2541 => x"74",
          2542 => x"0c",
          2543 => x"04",
          2544 => x"66",
          2545 => x"78",
          2546 => x"5a",
          2547 => x"80",
          2548 => x"38",
          2549 => x"09",
          2550 => x"e4",
          2551 => x"7a",
          2552 => x"5c",
          2553 => x"5b",
          2554 => x"09",
          2555 => x"38",
          2556 => x"39",
          2557 => x"09",
          2558 => x"38",
          2559 => x"70",
          2560 => x"33",
          2561 => x"2e",
          2562 => x"92",
          2563 => x"19",
          2564 => x"70",
          2565 => x"33",
          2566 => x"53",
          2567 => x"16",
          2568 => x"26",
          2569 => x"83",
          2570 => x"7c",
          2571 => x"05",
          2572 => x"05",
          2573 => x"5d",
          2574 => x"39",
          2575 => x"32",
          2576 => x"05",
          2577 => x"80",
          2578 => x"cc",
          2579 => x"81",
          2580 => x"07",
          2581 => x"07",
          2582 => x"51",
          2583 => x"80",
          2584 => x"79",
          2585 => x"70",
          2586 => x"33",
          2587 => x"80",
          2588 => x"38",
          2589 => x"e0",
          2590 => x"38",
          2591 => x"81",
          2592 => x"53",
          2593 => x"2e",
          2594 => x"73",
          2595 => x"a2",
          2596 => x"c3",
          2597 => x"38",
          2598 => x"24",
          2599 => x"80",
          2600 => x"8c",
          2601 => x"39",
          2602 => x"2e",
          2603 => x"81",
          2604 => x"80",
          2605 => x"80",
          2606 => x"d5",
          2607 => x"73",
          2608 => x"8e",
          2609 => x"39",
          2610 => x"2e",
          2611 => x"80",
          2612 => x"84",
          2613 => x"56",
          2614 => x"74",
          2615 => x"72",
          2616 => x"38",
          2617 => x"15",
          2618 => x"54",
          2619 => x"38",
          2620 => x"56",
          2621 => x"81",
          2622 => x"72",
          2623 => x"38",
          2624 => x"8a",
          2625 => x"06",
          2626 => x"2e",
          2627 => x"51",
          2628 => x"74",
          2629 => x"53",
          2630 => x"fd",
          2631 => x"51",
          2632 => x"ef",
          2633 => x"19",
          2634 => x"53",
          2635 => x"39",
          2636 => x"39",
          2637 => x"39",
          2638 => x"39",
          2639 => x"39",
          2640 => x"ca",
          2641 => x"39",
          2642 => x"70",
          2643 => x"53",
          2644 => x"88",
          2645 => x"19",
          2646 => x"39",
          2647 => x"54",
          2648 => x"74",
          2649 => x"70",
          2650 => x"70",
          2651 => x"25",
          2652 => x"55",
          2653 => x"8f",
          2654 => x"2e",
          2655 => x"09",
          2656 => x"90",
          2657 => x"80",
          2658 => x"5e",
          2659 => x"74",
          2660 => x"3f",
          2661 => x"08",
          2662 => x"7c",
          2663 => x"54",
          2664 => x"82",
          2665 => x"55",
          2666 => x"92",
          2667 => x"53",
          2668 => x"2e",
          2669 => x"14",
          2670 => x"ff",
          2671 => x"14",
          2672 => x"70",
          2673 => x"34",
          2674 => x"09",
          2675 => x"77",
          2676 => x"51",
          2677 => x"9f",
          2678 => x"72",
          2679 => x"79",
          2680 => x"81",
          2681 => x"72",
          2682 => x"38",
          2683 => x"05",
          2684 => x"ad",
          2685 => x"17",
          2686 => x"81",
          2687 => x"b0",
          2688 => x"38",
          2689 => x"81",
          2690 => x"06",
          2691 => x"9f",
          2692 => x"55",
          2693 => x"97",
          2694 => x"f9",
          2695 => x"81",
          2696 => x"8b",
          2697 => x"16",
          2698 => x"73",
          2699 => x"96",
          2700 => x"e0",
          2701 => x"17",
          2702 => x"33",
          2703 => x"f9",
          2704 => x"f2",
          2705 => x"16",
          2706 => x"7b",
          2707 => x"38",
          2708 => x"ba",
          2709 => x"96",
          2710 => x"fd",
          2711 => x"3d",
          2712 => x"05",
          2713 => x"52",
          2714 => x"d4",
          2715 => x"0d",
          2716 => x"0d",
          2717 => x"fc",
          2718 => x"88",
          2719 => x"51",
          2720 => x"82",
          2721 => x"53",
          2722 => x"80",
          2723 => x"fc",
          2724 => x"0d",
          2725 => x"0d",
          2726 => x"08",
          2727 => x"f4",
          2728 => x"88",
          2729 => x"52",
          2730 => x"3f",
          2731 => x"f4",
          2732 => x"0d",
          2733 => x"0d",
          2734 => x"9c",
          2735 => x"56",
          2736 => x"80",
          2737 => x"2e",
          2738 => x"82",
          2739 => x"52",
          2740 => x"85",
          2741 => x"ff",
          2742 => x"80",
          2743 => x"38",
          2744 => x"bc",
          2745 => x"32",
          2746 => x"05",
          2747 => x"51",
          2748 => x"80",
          2749 => x"71",
          2750 => x"38",
          2751 => x"98",
          2752 => x"25",
          2753 => x"16",
          2754 => x"25",
          2755 => x"74",
          2756 => x"72",
          2757 => x"54",
          2758 => x"f2",
          2759 => x"39",
          2760 => x"80",
          2761 => x"51",
          2762 => x"81",
          2763 => x"85",
          2764 => x"3d",
          2765 => x"3d",
          2766 => x"f8",
          2767 => x"9c",
          2768 => x"53",
          2769 => x"fe",
          2770 => x"82",
          2771 => x"84",
          2772 => x"f8",
          2773 => x"7c",
          2774 => x"70",
          2775 => x"75",
          2776 => x"55",
          2777 => x"2e",
          2778 => x"87",
          2779 => x"76",
          2780 => x"73",
          2781 => x"81",
          2782 => x"81",
          2783 => x"77",
          2784 => x"70",
          2785 => x"58",
          2786 => x"09",
          2787 => x"c2",
          2788 => x"81",
          2789 => x"75",
          2790 => x"55",
          2791 => x"e2",
          2792 => x"90",
          2793 => x"f8",
          2794 => x"8f",
          2795 => x"81",
          2796 => x"75",
          2797 => x"55",
          2798 => x"81",
          2799 => x"27",
          2800 => x"d0",
          2801 => x"55",
          2802 => x"73",
          2803 => x"80",
          2804 => x"14",
          2805 => x"72",
          2806 => x"ea",
          2807 => x"80",
          2808 => x"39",
          2809 => x"55",
          2810 => x"80",
          2811 => x"e0",
          2812 => x"38",
          2813 => x"81",
          2814 => x"53",
          2815 => x"81",
          2816 => x"53",
          2817 => x"8e",
          2818 => x"70",
          2819 => x"55",
          2820 => x"27",
          2821 => x"77",
          2822 => x"76",
          2823 => x"c4",
          2824 => x"85",
          2825 => x"76",
          2826 => x"77",
          2827 => x"70",
          2828 => x"55",
          2829 => x"77",
          2830 => x"38",
          2831 => x"05",
          2832 => x"0c",
          2833 => x"82",
          2834 => x"8a",
          2835 => x"f8",
          2836 => x"7c",
          2837 => x"70",
          2838 => x"75",
          2839 => x"55",
          2840 => x"2e",
          2841 => x"87",
          2842 => x"76",
          2843 => x"73",
          2844 => x"81",
          2845 => x"81",
          2846 => x"77",
          2847 => x"70",
          2848 => x"58",
          2849 => x"09",
          2850 => x"c2",
          2851 => x"81",
          2852 => x"75",
          2853 => x"55",
          2854 => x"e2",
          2855 => x"90",
          2856 => x"f8",
          2857 => x"8f",
          2858 => x"81",
          2859 => x"75",
          2860 => x"55",
          2861 => x"81",
          2862 => x"27",
          2863 => x"d0",
          2864 => x"55",
          2865 => x"73",
          2866 => x"80",
          2867 => x"14",
          2868 => x"72",
          2869 => x"ea",
          2870 => x"80",
          2871 => x"39",
          2872 => x"55",
          2873 => x"80",
          2874 => x"e0",
          2875 => x"38",
          2876 => x"81",
          2877 => x"53",
          2878 => x"81",
          2879 => x"53",
          2880 => x"8e",
          2881 => x"70",
          2882 => x"55",
          2883 => x"27",
          2884 => x"77",
          2885 => x"76",
          2886 => x"c2",
          2887 => x"85",
          2888 => x"76",
          2889 => x"77",
          2890 => x"70",
          2891 => x"55",
          2892 => x"77",
          2893 => x"38",
          2894 => x"05",
          2895 => x"0c",
          2896 => x"82",
          2897 => x"8a",
          2898 => x"fd",
          2899 => x"98",
          2900 => x"2c",
          2901 => x"70",
          2902 => x"10",
          2903 => x"2b",
          2904 => x"55",
          2905 => x"0b",
          2906 => x"12",
          2907 => x"72",
          2908 => x"38",
          2909 => x"f4",
          2910 => x"02",
          2911 => x"05",
          2912 => x"52",
          2913 => x"70",
          2914 => x"81",
          2915 => x"81",
          2916 => x"71",
          2917 => x"0c",
          2918 => x"04",
          2919 => x"78",
          2920 => x"9f",
          2921 => x"33",
          2922 => x"71",
          2923 => x"38",
          2924 => x"da",
          2925 => x"f2",
          2926 => x"51",
          2927 => x"72",
          2928 => x"52",
          2929 => x"71",
          2930 => x"52",
          2931 => x"51",
          2932 => x"73",
          2933 => x"3d",
          2934 => x"3d",
          2935 => x"84",
          2936 => x"33",
          2937 => x"bb",
          2938 => x"85",
          2939 => x"82",
          2940 => x"ec",
          2941 => x"59",
          2942 => x"59",
          2943 => x"86",
          2944 => x"9a",
          2945 => x"85",
          2946 => x"82",
          2947 => x"ec",
          2948 => x"70",
          2949 => x"56",
          2950 => x"3f",
          2951 => x"08",
          2952 => x"85",
          2953 => x"82",
          2954 => x"ec",
          2955 => x"56",
          2956 => x"2e",
          2957 => x"53",
          2958 => x"51",
          2959 => x"3f",
          2960 => x"33",
          2961 => x"74",
          2962 => x"34",
          2963 => x"06",
          2964 => x"27",
          2965 => x"0b",
          2966 => x"34",
          2967 => x"b6",
          2968 => x"c0",
          2969 => x"80",
          2970 => x"82",
          2971 => x"55",
          2972 => x"8c",
          2973 => x"54",
          2974 => x"52",
          2975 => x"d5",
          2976 => x"85",
          2977 => x"8a",
          2978 => x"cd",
          2979 => x"c0",
          2980 => x"d8",
          2981 => x"3d",
          2982 => x"3d",
          2983 => x"ec",
          2984 => x"72",
          2985 => x"80",
          2986 => x"71",
          2987 => x"3f",
          2988 => x"ff",
          2989 => x"54",
          2990 => x"25",
          2991 => x"0b",
          2992 => x"34",
          2993 => x"08",
          2994 => x"2e",
          2995 => x"51",
          2996 => x"3f",
          2997 => x"08",
          2998 => x"3f",
          2999 => x"85",
          3000 => x"3d",
          3001 => x"3d",
          3002 => x"80",
          3003 => x"c0",
          3004 => x"de",
          3005 => x"85",
          3006 => x"d2",
          3007 => x"c0",
          3008 => x"f8",
          3009 => x"70",
          3010 => x"87",
          3011 => x"85",
          3012 => x"2e",
          3013 => x"51",
          3014 => x"3f",
          3015 => x"08",
          3016 => x"82",
          3017 => x"25",
          3018 => x"85",
          3019 => x"05",
          3020 => x"55",
          3021 => x"75",
          3022 => x"81",
          3023 => x"e8",
          3024 => x"97",
          3025 => x"2e",
          3026 => x"ff",
          3027 => x"3d",
          3028 => x"3d",
          3029 => x"08",
          3030 => x"5a",
          3031 => x"58",
          3032 => x"82",
          3033 => x"51",
          3034 => x"3f",
          3035 => x"08",
          3036 => x"ff",
          3037 => x"c0",
          3038 => x"80",
          3039 => x"3d",
          3040 => x"81",
          3041 => x"82",
          3042 => x"80",
          3043 => x"75",
          3044 => x"a5",
          3045 => x"ec",
          3046 => x"58",
          3047 => x"82",
          3048 => x"25",
          3049 => x"85",
          3050 => x"05",
          3051 => x"55",
          3052 => x"74",
          3053 => x"81",
          3054 => x"07",
          3055 => x"55",
          3056 => x"2e",
          3057 => x"ff",
          3058 => x"85",
          3059 => x"11",
          3060 => x"80",
          3061 => x"82",
          3062 => x"80",
          3063 => x"81",
          3064 => x"ef",
          3065 => x"77",
          3066 => x"06",
          3067 => x"52",
          3068 => x"b4",
          3069 => x"51",
          3070 => x"3f",
          3071 => x"54",
          3072 => x"08",
          3073 => x"58",
          3074 => x"ec",
          3075 => x"0d",
          3076 => x"0d",
          3077 => x"5c",
          3078 => x"57",
          3079 => x"73",
          3080 => x"81",
          3081 => x"78",
          3082 => x"56",
          3083 => x"98",
          3084 => x"70",
          3085 => x"33",
          3086 => x"73",
          3087 => x"81",
          3088 => x"75",
          3089 => x"38",
          3090 => x"83",
          3091 => x"c8",
          3092 => x"53",
          3093 => x"b2",
          3094 => x"85",
          3095 => x"79",
          3096 => x"51",
          3097 => x"3f",
          3098 => x"08",
          3099 => x"84",
          3100 => x"73",
          3101 => x"38",
          3102 => x"88",
          3103 => x"fc",
          3104 => x"39",
          3105 => x"8c",
          3106 => x"53",
          3107 => x"f5",
          3108 => x"85",
          3109 => x"2e",
          3110 => x"1b",
          3111 => x"77",
          3112 => x"3f",
          3113 => x"08",
          3114 => x"54",
          3115 => x"91",
          3116 => x"70",
          3117 => x"56",
          3118 => x"27",
          3119 => x"80",
          3120 => x"85",
          3121 => x"3d",
          3122 => x"3d",
          3123 => x"08",
          3124 => x"b4",
          3125 => x"5f",
          3126 => x"af",
          3127 => x"85",
          3128 => x"85",
          3129 => x"5b",
          3130 => x"38",
          3131 => x"bc",
          3132 => x"73",
          3133 => x"55",
          3134 => x"81",
          3135 => x"70",
          3136 => x"56",
          3137 => x"81",
          3138 => x"51",
          3139 => x"82",
          3140 => x"82",
          3141 => x"82",
          3142 => x"80",
          3143 => x"38",
          3144 => x"52",
          3145 => x"08",
          3146 => x"90",
          3147 => x"ec",
          3148 => x"8b",
          3149 => x"a0",
          3150 => x"3f",
          3151 => x"82",
          3152 => x"5b",
          3153 => x"08",
          3154 => x"52",
          3155 => x"52",
          3156 => x"ec",
          3157 => x"ec",
          3158 => x"85",
          3159 => x"2e",
          3160 => x"80",
          3161 => x"85",
          3162 => x"ff",
          3163 => x"82",
          3164 => x"55",
          3165 => x"85",
          3166 => x"a9",
          3167 => x"ec",
          3168 => x"70",
          3169 => x"80",
          3170 => x"53",
          3171 => x"06",
          3172 => x"f8",
          3173 => x"1b",
          3174 => x"06",
          3175 => x"7b",
          3176 => x"80",
          3177 => x"2e",
          3178 => x"ff",
          3179 => x"39",
          3180 => x"bc",
          3181 => x"38",
          3182 => x"08",
          3183 => x"38",
          3184 => x"8f",
          3185 => x"9c",
          3186 => x"ec",
          3187 => x"70",
          3188 => x"59",
          3189 => x"ee",
          3190 => x"ff",
          3191 => x"84",
          3192 => x"2b",
          3193 => x"82",
          3194 => x"70",
          3195 => x"97",
          3196 => x"2c",
          3197 => x"2b",
          3198 => x"11",
          3199 => x"33",
          3200 => x"51",
          3201 => x"59",
          3202 => x"56",
          3203 => x"80",
          3204 => x"74",
          3205 => x"ff",
          3206 => x"2b",
          3207 => x"51",
          3208 => x"75",
          3209 => x"38",
          3210 => x"52",
          3211 => x"9b",
          3212 => x"ec",
          3213 => x"06",
          3214 => x"2e",
          3215 => x"82",
          3216 => x"81",
          3217 => x"81",
          3218 => x"2b",
          3219 => x"70",
          3220 => x"53",
          3221 => x"73",
          3222 => x"38",
          3223 => x"52",
          3224 => x"e7",
          3225 => x"ec",
          3226 => x"06",
          3227 => x"38",
          3228 => x"56",
          3229 => x"80",
          3230 => x"1c",
          3231 => x"9d",
          3232 => x"98",
          3233 => x"2c",
          3234 => x"33",
          3235 => x"70",
          3236 => x"10",
          3237 => x"2b",
          3238 => x"11",
          3239 => x"53",
          3240 => x"51",
          3241 => x"2e",
          3242 => x"fe",
          3243 => x"fa",
          3244 => x"7d",
          3245 => x"82",
          3246 => x"80",
          3247 => x"80",
          3248 => x"75",
          3249 => x"34",
          3250 => x"80",
          3251 => x"3d",
          3252 => x"0c",
          3253 => x"95",
          3254 => x"38",
          3255 => x"54",
          3256 => x"14",
          3257 => x"9d",
          3258 => x"75",
          3259 => x"d3",
          3260 => x"88",
          3261 => x"74",
          3262 => x"73",
          3263 => x"98",
          3264 => x"75",
          3265 => x"38",
          3266 => x"73",
          3267 => x"34",
          3268 => x"98",
          3269 => x"2c",
          3270 => x"33",
          3271 => x"54",
          3272 => x"e4",
          3273 => x"8c",
          3274 => x"56",
          3275 => x"9d",
          3276 => x"1a",
          3277 => x"33",
          3278 => x"9d",
          3279 => x"73",
          3280 => x"38",
          3281 => x"73",
          3282 => x"34",
          3283 => x"33",
          3284 => x"98",
          3285 => x"2c",
          3286 => x"33",
          3287 => x"54",
          3288 => x"9f",
          3289 => x"70",
          3290 => x"e7",
          3291 => x"15",
          3292 => x"70",
          3293 => x"9d",
          3294 => x"51",
          3295 => x"75",
          3296 => x"82",
          3297 => x"70",
          3298 => x"98",
          3299 => x"88",
          3300 => x"56",
          3301 => x"25",
          3302 => x"88",
          3303 => x"3f",
          3304 => x"98",
          3305 => x"2c",
          3306 => x"33",
          3307 => x"54",
          3308 => x"e7",
          3309 => x"39",
          3310 => x"80",
          3311 => x"34",
          3312 => x"53",
          3313 => x"f3",
          3314 => x"d0",
          3315 => x"39",
          3316 => x"33",
          3317 => x"06",
          3318 => x"80",
          3319 => x"38",
          3320 => x"33",
          3321 => x"73",
          3322 => x"34",
          3323 => x"73",
          3324 => x"34",
          3325 => x"96",
          3326 => x"8c",
          3327 => x"2b",
          3328 => x"82",
          3329 => x"57",
          3330 => x"74",
          3331 => x"38",
          3332 => x"81",
          3333 => x"34",
          3334 => x"e5",
          3335 => x"15",
          3336 => x"70",
          3337 => x"9d",
          3338 => x"51",
          3339 => x"75",
          3340 => x"a0",
          3341 => x"3f",
          3342 => x"33",
          3343 => x"70",
          3344 => x"9d",
          3345 => x"51",
          3346 => x"74",
          3347 => x"38",
          3348 => x"ba",
          3349 => x"70",
          3350 => x"98",
          3351 => x"88",
          3352 => x"56",
          3353 => x"25",
          3354 => x"d7",
          3355 => x"88",
          3356 => x"54",
          3357 => x"8a",
          3358 => x"3f",
          3359 => x"52",
          3360 => x"8d",
          3361 => x"ec",
          3362 => x"06",
          3363 => x"38",
          3364 => x"33",
          3365 => x"2e",
          3366 => x"53",
          3367 => x"51",
          3368 => x"84",
          3369 => x"34",
          3370 => x"9d",
          3371 => x"0b",
          3372 => x"34",
          3373 => x"ec",
          3374 => x"0d",
          3375 => x"8c",
          3376 => x"80",
          3377 => x"38",
          3378 => x"c2",
          3379 => x"8c",
          3380 => x"54",
          3381 => x"8c",
          3382 => x"ff",
          3383 => x"39",
          3384 => x"33",
          3385 => x"33",
          3386 => x"75",
          3387 => x"38",
          3388 => x"73",
          3389 => x"34",
          3390 => x"70",
          3391 => x"81",
          3392 => x"51",
          3393 => x"25",
          3394 => x"1a",
          3395 => x"33",
          3396 => x"33",
          3397 => x"3f",
          3398 => x"98",
          3399 => x"2c",
          3400 => x"33",
          3401 => x"54",
          3402 => x"de",
          3403 => x"e3",
          3404 => x"9d",
          3405 => x"98",
          3406 => x"2c",
          3407 => x"33",
          3408 => x"57",
          3409 => x"f8",
          3410 => x"51",
          3411 => x"81",
          3412 => x"2b",
          3413 => x"82",
          3414 => x"59",
          3415 => x"75",
          3416 => x"38",
          3417 => x"82",
          3418 => x"70",
          3419 => x"82",
          3420 => x"59",
          3421 => x"77",
          3422 => x"38",
          3423 => x"73",
          3424 => x"34",
          3425 => x"33",
          3426 => x"82",
          3427 => x"8c",
          3428 => x"ff",
          3429 => x"88",
          3430 => x"54",
          3431 => x"dc",
          3432 => x"39",
          3433 => x"53",
          3434 => x"f3",
          3435 => x"ec",
          3436 => x"82",
          3437 => x"80",
          3438 => x"88",
          3439 => x"39",
          3440 => x"82",
          3441 => x"55",
          3442 => x"a6",
          3443 => x"ff",
          3444 => x"82",
          3445 => x"82",
          3446 => x"82",
          3447 => x"81",
          3448 => x"05",
          3449 => x"79",
          3450 => x"ad",
          3451 => x"81",
          3452 => x"82",
          3453 => x"ec",
          3454 => x"08",
          3455 => x"74",
          3456 => x"38",
          3457 => x"a7",
          3458 => x"85",
          3459 => x"9d",
          3460 => x"85",
          3461 => x"ff",
          3462 => x"53",
          3463 => x"51",
          3464 => x"3f",
          3465 => x"80",
          3466 => x"08",
          3467 => x"2e",
          3468 => x"74",
          3469 => x"81",
          3470 => x"7a",
          3471 => x"81",
          3472 => x"82",
          3473 => x"55",
          3474 => x"a4",
          3475 => x"ff",
          3476 => x"82",
          3477 => x"82",
          3478 => x"82",
          3479 => x"81",
          3480 => x"05",
          3481 => x"79",
          3482 => x"ad",
          3483 => x"39",
          3484 => x"82",
          3485 => x"08",
          3486 => x"80",
          3487 => x"74",
          3488 => x"b5",
          3489 => x"ec",
          3490 => x"88",
          3491 => x"ec",
          3492 => x"06",
          3493 => x"74",
          3494 => x"ff",
          3495 => x"81",
          3496 => x"81",
          3497 => x"89",
          3498 => x"9d",
          3499 => x"7a",
          3500 => x"8c",
          3501 => x"88",
          3502 => x"51",
          3503 => x"f6",
          3504 => x"9d",
          3505 => x"81",
          3506 => x"9d",
          3507 => x"56",
          3508 => x"27",
          3509 => x"81",
          3510 => x"82",
          3511 => x"74",
          3512 => x"52",
          3513 => x"3f",
          3514 => x"82",
          3515 => x"54",
          3516 => x"f5",
          3517 => x"51",
          3518 => x"82",
          3519 => x"ff",
          3520 => x"82",
          3521 => x"f5",
          3522 => x"3d",
          3523 => x"f4",
          3524 => x"e4",
          3525 => x"0b",
          3526 => x"23",
          3527 => x"80",
          3528 => x"f4",
          3529 => x"c5",
          3530 => x"e4",
          3531 => x"58",
          3532 => x"81",
          3533 => x"15",
          3534 => x"e4",
          3535 => x"84",
          3536 => x"85",
          3537 => x"85",
          3538 => x"77",
          3539 => x"76",
          3540 => x"82",
          3541 => x"82",
          3542 => x"ff",
          3543 => x"80",
          3544 => x"ff",
          3545 => x"88",
          3546 => x"55",
          3547 => x"17",
          3548 => x"17",
          3549 => x"e0",
          3550 => x"2b",
          3551 => x"08",
          3552 => x"51",
          3553 => x"82",
          3554 => x"83",
          3555 => x"3d",
          3556 => x"3d",
          3557 => x"81",
          3558 => x"27",
          3559 => x"12",
          3560 => x"11",
          3561 => x"ff",
          3562 => x"51",
          3563 => x"ec",
          3564 => x"0d",
          3565 => x"0d",
          3566 => x"22",
          3567 => x"aa",
          3568 => x"05",
          3569 => x"08",
          3570 => x"71",
          3571 => x"2b",
          3572 => x"33",
          3573 => x"71",
          3574 => x"02",
          3575 => x"05",
          3576 => x"ff",
          3577 => x"70",
          3578 => x"51",
          3579 => x"5b",
          3580 => x"54",
          3581 => x"34",
          3582 => x"34",
          3583 => x"08",
          3584 => x"2a",
          3585 => x"82",
          3586 => x"83",
          3587 => x"85",
          3588 => x"17",
          3589 => x"12",
          3590 => x"2b",
          3591 => x"2b",
          3592 => x"06",
          3593 => x"52",
          3594 => x"83",
          3595 => x"70",
          3596 => x"54",
          3597 => x"12",
          3598 => x"ff",
          3599 => x"83",
          3600 => x"85",
          3601 => x"56",
          3602 => x"72",
          3603 => x"89",
          3604 => x"fb",
          3605 => x"85",
          3606 => x"84",
          3607 => x"22",
          3608 => x"72",
          3609 => x"33",
          3610 => x"71",
          3611 => x"83",
          3612 => x"5b",
          3613 => x"52",
          3614 => x"12",
          3615 => x"33",
          3616 => x"07",
          3617 => x"54",
          3618 => x"70",
          3619 => x"73",
          3620 => x"82",
          3621 => x"70",
          3622 => x"33",
          3623 => x"71",
          3624 => x"83",
          3625 => x"59",
          3626 => x"05",
          3627 => x"87",
          3628 => x"88",
          3629 => x"88",
          3630 => x"56",
          3631 => x"13",
          3632 => x"13",
          3633 => x"e4",
          3634 => x"33",
          3635 => x"71",
          3636 => x"70",
          3637 => x"06",
          3638 => x"53",
          3639 => x"53",
          3640 => x"70",
          3641 => x"87",
          3642 => x"f9",
          3643 => x"a6",
          3644 => x"85",
          3645 => x"83",
          3646 => x"70",
          3647 => x"33",
          3648 => x"07",
          3649 => x"53",
          3650 => x"58",
          3651 => x"33",
          3652 => x"71",
          3653 => x"90",
          3654 => x"5a",
          3655 => x"71",
          3656 => x"f6",
          3657 => x"fe",
          3658 => x"85",
          3659 => x"17",
          3660 => x"12",
          3661 => x"2b",
          3662 => x"07",
          3663 => x"33",
          3664 => x"71",
          3665 => x"70",
          3666 => x"ff",
          3667 => x"52",
          3668 => x"57",
          3669 => x"05",
          3670 => x"54",
          3671 => x"13",
          3672 => x"13",
          3673 => x"e4",
          3674 => x"70",
          3675 => x"33",
          3676 => x"71",
          3677 => x"56",
          3678 => x"72",
          3679 => x"81",
          3680 => x"88",
          3681 => x"81",
          3682 => x"70",
          3683 => x"51",
          3684 => x"72",
          3685 => x"81",
          3686 => x"3d",
          3687 => x"3d",
          3688 => x"e4",
          3689 => x"05",
          3690 => x"70",
          3691 => x"11",
          3692 => x"83",
          3693 => x"8b",
          3694 => x"2b",
          3695 => x"59",
          3696 => x"73",
          3697 => x"81",
          3698 => x"88",
          3699 => x"8c",
          3700 => x"22",
          3701 => x"88",
          3702 => x"53",
          3703 => x"73",
          3704 => x"14",
          3705 => x"e4",
          3706 => x"70",
          3707 => x"33",
          3708 => x"71",
          3709 => x"56",
          3710 => x"72",
          3711 => x"33",
          3712 => x"71",
          3713 => x"70",
          3714 => x"55",
          3715 => x"82",
          3716 => x"83",
          3717 => x"85",
          3718 => x"82",
          3719 => x"12",
          3720 => x"2b",
          3721 => x"ec",
          3722 => x"87",
          3723 => x"f7",
          3724 => x"82",
          3725 => x"31",
          3726 => x"83",
          3727 => x"70",
          3728 => x"fd",
          3729 => x"85",
          3730 => x"83",
          3731 => x"82",
          3732 => x"12",
          3733 => x"2b",
          3734 => x"07",
          3735 => x"33",
          3736 => x"71",
          3737 => x"90",
          3738 => x"42",
          3739 => x"5b",
          3740 => x"54",
          3741 => x"8d",
          3742 => x"80",
          3743 => x"fe",
          3744 => x"84",
          3745 => x"33",
          3746 => x"71",
          3747 => x"83",
          3748 => x"11",
          3749 => x"53",
          3750 => x"55",
          3751 => x"34",
          3752 => x"06",
          3753 => x"14",
          3754 => x"e4",
          3755 => x"84",
          3756 => x"13",
          3757 => x"2b",
          3758 => x"2a",
          3759 => x"56",
          3760 => x"16",
          3761 => x"16",
          3762 => x"e4",
          3763 => x"80",
          3764 => x"34",
          3765 => x"14",
          3766 => x"e4",
          3767 => x"84",
          3768 => x"85",
          3769 => x"85",
          3770 => x"70",
          3771 => x"33",
          3772 => x"07",
          3773 => x"80",
          3774 => x"2a",
          3775 => x"56",
          3776 => x"34",
          3777 => x"34",
          3778 => x"04",
          3779 => x"73",
          3780 => x"e4",
          3781 => x"f7",
          3782 => x"80",
          3783 => x"71",
          3784 => x"3f",
          3785 => x"04",
          3786 => x"80",
          3787 => x"f8",
          3788 => x"85",
          3789 => x"ff",
          3790 => x"85",
          3791 => x"11",
          3792 => x"33",
          3793 => x"07",
          3794 => x"56",
          3795 => x"ff",
          3796 => x"78",
          3797 => x"38",
          3798 => x"77",
          3799 => x"81",
          3800 => x"88",
          3801 => x"81",
          3802 => x"79",
          3803 => x"ff",
          3804 => x"7f",
          3805 => x"51",
          3806 => x"77",
          3807 => x"38",
          3808 => x"85",
          3809 => x"5a",
          3810 => x"33",
          3811 => x"71",
          3812 => x"57",
          3813 => x"38",
          3814 => x"ff",
          3815 => x"7a",
          3816 => x"80",
          3817 => x"82",
          3818 => x"11",
          3819 => x"12",
          3820 => x"2b",
          3821 => x"ff",
          3822 => x"52",
          3823 => x"55",
          3824 => x"83",
          3825 => x"80",
          3826 => x"26",
          3827 => x"74",
          3828 => x"2e",
          3829 => x"77",
          3830 => x"81",
          3831 => x"75",
          3832 => x"3f",
          3833 => x"82",
          3834 => x"79",
          3835 => x"f7",
          3836 => x"85",
          3837 => x"1c",
          3838 => x"87",
          3839 => x"8b",
          3840 => x"2b",
          3841 => x"5e",
          3842 => x"7a",
          3843 => x"ff",
          3844 => x"88",
          3845 => x"56",
          3846 => x"15",
          3847 => x"ff",
          3848 => x"85",
          3849 => x"85",
          3850 => x"83",
          3851 => x"72",
          3852 => x"33",
          3853 => x"71",
          3854 => x"70",
          3855 => x"5b",
          3856 => x"56",
          3857 => x"19",
          3858 => x"19",
          3859 => x"e4",
          3860 => x"84",
          3861 => x"12",
          3862 => x"2b",
          3863 => x"07",
          3864 => x"55",
          3865 => x"78",
          3866 => x"76",
          3867 => x"82",
          3868 => x"70",
          3869 => x"84",
          3870 => x"12",
          3871 => x"2b",
          3872 => x"2a",
          3873 => x"52",
          3874 => x"84",
          3875 => x"85",
          3876 => x"85",
          3877 => x"84",
          3878 => x"82",
          3879 => x"8d",
          3880 => x"fe",
          3881 => x"52",
          3882 => x"08",
          3883 => x"da",
          3884 => x"71",
          3885 => x"38",
          3886 => x"ec",
          3887 => x"ec",
          3888 => x"82",
          3889 => x"84",
          3890 => x"ff",
          3891 => x"8f",
          3892 => x"81",
          3893 => x"26",
          3894 => x"85",
          3895 => x"52",
          3896 => x"ec",
          3897 => x"0d",
          3898 => x"0d",
          3899 => x"33",
          3900 => x"9f",
          3901 => x"53",
          3902 => x"81",
          3903 => x"38",
          3904 => x"87",
          3905 => x"11",
          3906 => x"54",
          3907 => x"84",
          3908 => x"54",
          3909 => x"87",
          3910 => x"11",
          3911 => x"0c",
          3912 => x"c0",
          3913 => x"70",
          3914 => x"70",
          3915 => x"51",
          3916 => x"8a",
          3917 => x"98",
          3918 => x"70",
          3919 => x"08",
          3920 => x"06",
          3921 => x"38",
          3922 => x"8c",
          3923 => x"80",
          3924 => x"71",
          3925 => x"14",
          3926 => x"e8",
          3927 => x"70",
          3928 => x"0c",
          3929 => x"04",
          3930 => x"60",
          3931 => x"8c",
          3932 => x"33",
          3933 => x"5b",
          3934 => x"5a",
          3935 => x"82",
          3936 => x"81",
          3937 => x"52",
          3938 => x"38",
          3939 => x"84",
          3940 => x"92",
          3941 => x"c0",
          3942 => x"87",
          3943 => x"13",
          3944 => x"57",
          3945 => x"0b",
          3946 => x"8c",
          3947 => x"0c",
          3948 => x"75",
          3949 => x"2a",
          3950 => x"51",
          3951 => x"80",
          3952 => x"7b",
          3953 => x"7b",
          3954 => x"5d",
          3955 => x"59",
          3956 => x"06",
          3957 => x"73",
          3958 => x"81",
          3959 => x"ff",
          3960 => x"72",
          3961 => x"38",
          3962 => x"8c",
          3963 => x"c3",
          3964 => x"98",
          3965 => x"71",
          3966 => x"38",
          3967 => x"2e",
          3968 => x"76",
          3969 => x"92",
          3970 => x"72",
          3971 => x"06",
          3972 => x"f7",
          3973 => x"5a",
          3974 => x"80",
          3975 => x"70",
          3976 => x"5a",
          3977 => x"80",
          3978 => x"73",
          3979 => x"06",
          3980 => x"38",
          3981 => x"fe",
          3982 => x"fc",
          3983 => x"52",
          3984 => x"83",
          3985 => x"71",
          3986 => x"85",
          3987 => x"3d",
          3988 => x"3d",
          3989 => x"64",
          3990 => x"bf",
          3991 => x"40",
          3992 => x"59",
          3993 => x"58",
          3994 => x"82",
          3995 => x"81",
          3996 => x"52",
          3997 => x"09",
          3998 => x"b1",
          3999 => x"84",
          4000 => x"92",
          4001 => x"c0",
          4002 => x"87",
          4003 => x"13",
          4004 => x"56",
          4005 => x"87",
          4006 => x"0c",
          4007 => x"82",
          4008 => x"58",
          4009 => x"84",
          4010 => x"06",
          4011 => x"71",
          4012 => x"38",
          4013 => x"05",
          4014 => x"0c",
          4015 => x"73",
          4016 => x"81",
          4017 => x"71",
          4018 => x"38",
          4019 => x"8c",
          4020 => x"d0",
          4021 => x"98",
          4022 => x"71",
          4023 => x"38",
          4024 => x"2e",
          4025 => x"76",
          4026 => x"92",
          4027 => x"72",
          4028 => x"06",
          4029 => x"f7",
          4030 => x"59",
          4031 => x"1a",
          4032 => x"06",
          4033 => x"59",
          4034 => x"80",
          4035 => x"73",
          4036 => x"06",
          4037 => x"38",
          4038 => x"fe",
          4039 => x"fc",
          4040 => x"52",
          4041 => x"83",
          4042 => x"71",
          4043 => x"85",
          4044 => x"3d",
          4045 => x"3d",
          4046 => x"84",
          4047 => x"33",
          4048 => x"a7",
          4049 => x"54",
          4050 => x"fa",
          4051 => x"85",
          4052 => x"06",
          4053 => x"72",
          4054 => x"85",
          4055 => x"98",
          4056 => x"56",
          4057 => x"80",
          4058 => x"76",
          4059 => x"74",
          4060 => x"c0",
          4061 => x"54",
          4062 => x"2e",
          4063 => x"d4",
          4064 => x"2e",
          4065 => x"80",
          4066 => x"08",
          4067 => x"70",
          4068 => x"51",
          4069 => x"2e",
          4070 => x"c0",
          4071 => x"52",
          4072 => x"87",
          4073 => x"08",
          4074 => x"38",
          4075 => x"87",
          4076 => x"14",
          4077 => x"70",
          4078 => x"52",
          4079 => x"96",
          4080 => x"92",
          4081 => x"0a",
          4082 => x"39",
          4083 => x"0c",
          4084 => x"39",
          4085 => x"54",
          4086 => x"ec",
          4087 => x"0d",
          4088 => x"0d",
          4089 => x"33",
          4090 => x"88",
          4091 => x"85",
          4092 => x"51",
          4093 => x"04",
          4094 => x"75",
          4095 => x"82",
          4096 => x"90",
          4097 => x"2b",
          4098 => x"33",
          4099 => x"88",
          4100 => x"71",
          4101 => x"ec",
          4102 => x"54",
          4103 => x"85",
          4104 => x"ff",
          4105 => x"02",
          4106 => x"05",
          4107 => x"70",
          4108 => x"05",
          4109 => x"88",
          4110 => x"72",
          4111 => x"0d",
          4112 => x"0d",
          4113 => x"52",
          4114 => x"81",
          4115 => x"70",
          4116 => x"70",
          4117 => x"05",
          4118 => x"88",
          4119 => x"72",
          4120 => x"54",
          4121 => x"2a",
          4122 => x"34",
          4123 => x"04",
          4124 => x"76",
          4125 => x"54",
          4126 => x"2e",
          4127 => x"70",
          4128 => x"33",
          4129 => x"05",
          4130 => x"11",
          4131 => x"84",
          4132 => x"fe",
          4133 => x"77",
          4134 => x"53",
          4135 => x"81",
          4136 => x"ff",
          4137 => x"f4",
          4138 => x"0d",
          4139 => x"0d",
          4140 => x"56",
          4141 => x"70",
          4142 => x"33",
          4143 => x"05",
          4144 => x"71",
          4145 => x"56",
          4146 => x"72",
          4147 => x"38",
          4148 => x"e2",
          4149 => x"85",
          4150 => x"3d",
          4151 => x"3d",
          4152 => x"54",
          4153 => x"71",
          4154 => x"38",
          4155 => x"70",
          4156 => x"f3",
          4157 => x"82",
          4158 => x"84",
          4159 => x"80",
          4160 => x"ec",
          4161 => x"0b",
          4162 => x"0c",
          4163 => x"0d",
          4164 => x"0b",
          4165 => x"56",
          4166 => x"2e",
          4167 => x"81",
          4168 => x"08",
          4169 => x"70",
          4170 => x"33",
          4171 => x"a2",
          4172 => x"ec",
          4173 => x"09",
          4174 => x"38",
          4175 => x"08",
          4176 => x"b0",
          4177 => x"a4",
          4178 => x"9c",
          4179 => x"56",
          4180 => x"27",
          4181 => x"16",
          4182 => x"82",
          4183 => x"06",
          4184 => x"54",
          4185 => x"78",
          4186 => x"33",
          4187 => x"3f",
          4188 => x"5a",
          4189 => x"ec",
          4190 => x"0d",
          4191 => x"0d",
          4192 => x"56",
          4193 => x"b0",
          4194 => x"af",
          4195 => x"fe",
          4196 => x"85",
          4197 => x"82",
          4198 => x"9f",
          4199 => x"74",
          4200 => x"52",
          4201 => x"51",
          4202 => x"82",
          4203 => x"80",
          4204 => x"ff",
          4205 => x"74",
          4206 => x"76",
          4207 => x"0c",
          4208 => x"04",
          4209 => x"7a",
          4210 => x"fe",
          4211 => x"85",
          4212 => x"82",
          4213 => x"81",
          4214 => x"33",
          4215 => x"2e",
          4216 => x"80",
          4217 => x"17",
          4218 => x"81",
          4219 => x"06",
          4220 => x"84",
          4221 => x"85",
          4222 => x"b4",
          4223 => x"56",
          4224 => x"82",
          4225 => x"84",
          4226 => x"fc",
          4227 => x"8b",
          4228 => x"52",
          4229 => x"a9",
          4230 => x"85",
          4231 => x"84",
          4232 => x"fc",
          4233 => x"17",
          4234 => x"9c",
          4235 => x"91",
          4236 => x"08",
          4237 => x"17",
          4238 => x"3f",
          4239 => x"81",
          4240 => x"19",
          4241 => x"53",
          4242 => x"17",
          4243 => x"82",
          4244 => x"18",
          4245 => x"80",
          4246 => x"33",
          4247 => x"3f",
          4248 => x"08",
          4249 => x"38",
          4250 => x"82",
          4251 => x"8a",
          4252 => x"fb",
          4253 => x"fe",
          4254 => x"08",
          4255 => x"55",
          4256 => x"73",
          4257 => x"38",
          4258 => x"74",
          4259 => x"97",
          4260 => x"15",
          4261 => x"ec",
          4262 => x"75",
          4263 => x"0c",
          4264 => x"04",
          4265 => x"7a",
          4266 => x"56",
          4267 => x"77",
          4268 => x"38",
          4269 => x"08",
          4270 => x"38",
          4271 => x"54",
          4272 => x"2e",
          4273 => x"72",
          4274 => x"38",
          4275 => x"8d",
          4276 => x"39",
          4277 => x"81",
          4278 => x"b6",
          4279 => x"2a",
          4280 => x"2a",
          4281 => x"05",
          4282 => x"55",
          4283 => x"82",
          4284 => x"81",
          4285 => x"83",
          4286 => x"b4",
          4287 => x"17",
          4288 => x"a4",
          4289 => x"55",
          4290 => x"57",
          4291 => x"3f",
          4292 => x"08",
          4293 => x"74",
          4294 => x"14",
          4295 => x"70",
          4296 => x"07",
          4297 => x"71",
          4298 => x"52",
          4299 => x"72",
          4300 => x"75",
          4301 => x"58",
          4302 => x"76",
          4303 => x"15",
          4304 => x"73",
          4305 => x"3f",
          4306 => x"08",
          4307 => x"76",
          4308 => x"06",
          4309 => x"05",
          4310 => x"3f",
          4311 => x"08",
          4312 => x"06",
          4313 => x"76",
          4314 => x"15",
          4315 => x"73",
          4316 => x"3f",
          4317 => x"08",
          4318 => x"82",
          4319 => x"06",
          4320 => x"05",
          4321 => x"3f",
          4322 => x"08",
          4323 => x"58",
          4324 => x"58",
          4325 => x"ec",
          4326 => x"0d",
          4327 => x"0d",
          4328 => x"5a",
          4329 => x"59",
          4330 => x"82",
          4331 => x"98",
          4332 => x"82",
          4333 => x"33",
          4334 => x"2e",
          4335 => x"72",
          4336 => x"38",
          4337 => x"8d",
          4338 => x"39",
          4339 => x"81",
          4340 => x"f7",
          4341 => x"2a",
          4342 => x"2a",
          4343 => x"05",
          4344 => x"55",
          4345 => x"82",
          4346 => x"59",
          4347 => x"08",
          4348 => x"74",
          4349 => x"16",
          4350 => x"16",
          4351 => x"59",
          4352 => x"53",
          4353 => x"8f",
          4354 => x"2b",
          4355 => x"74",
          4356 => x"71",
          4357 => x"72",
          4358 => x"0b",
          4359 => x"74",
          4360 => x"17",
          4361 => x"75",
          4362 => x"3f",
          4363 => x"08",
          4364 => x"ec",
          4365 => x"38",
          4366 => x"06",
          4367 => x"78",
          4368 => x"54",
          4369 => x"77",
          4370 => x"33",
          4371 => x"71",
          4372 => x"51",
          4373 => x"34",
          4374 => x"76",
          4375 => x"17",
          4376 => x"75",
          4377 => x"3f",
          4378 => x"08",
          4379 => x"ec",
          4380 => x"38",
          4381 => x"ff",
          4382 => x"10",
          4383 => x"76",
          4384 => x"51",
          4385 => x"be",
          4386 => x"2a",
          4387 => x"05",
          4388 => x"f9",
          4389 => x"85",
          4390 => x"82",
          4391 => x"ab",
          4392 => x"0a",
          4393 => x"2b",
          4394 => x"70",
          4395 => x"70",
          4396 => x"54",
          4397 => x"82",
          4398 => x"8f",
          4399 => x"07",
          4400 => x"f6",
          4401 => x"0b",
          4402 => x"78",
          4403 => x"0c",
          4404 => x"04",
          4405 => x"7a",
          4406 => x"08",
          4407 => x"59",
          4408 => x"a4",
          4409 => x"17",
          4410 => x"38",
          4411 => x"aa",
          4412 => x"73",
          4413 => x"fd",
          4414 => x"85",
          4415 => x"82",
          4416 => x"80",
          4417 => x"39",
          4418 => x"eb",
          4419 => x"80",
          4420 => x"85",
          4421 => x"80",
          4422 => x"52",
          4423 => x"84",
          4424 => x"ec",
          4425 => x"85",
          4426 => x"2e",
          4427 => x"82",
          4428 => x"81",
          4429 => x"82",
          4430 => x"ff",
          4431 => x"80",
          4432 => x"75",
          4433 => x"3f",
          4434 => x"08",
          4435 => x"16",
          4436 => x"90",
          4437 => x"55",
          4438 => x"27",
          4439 => x"15",
          4440 => x"84",
          4441 => x"07",
          4442 => x"17",
          4443 => x"76",
          4444 => x"a6",
          4445 => x"73",
          4446 => x"0c",
          4447 => x"04",
          4448 => x"7c",
          4449 => x"59",
          4450 => x"95",
          4451 => x"08",
          4452 => x"2e",
          4453 => x"17",
          4454 => x"b2",
          4455 => x"ae",
          4456 => x"7a",
          4457 => x"3f",
          4458 => x"82",
          4459 => x"27",
          4460 => x"82",
          4461 => x"55",
          4462 => x"08",
          4463 => x"d8",
          4464 => x"08",
          4465 => x"08",
          4466 => x"38",
          4467 => x"17",
          4468 => x"54",
          4469 => x"82",
          4470 => x"7a",
          4471 => x"06",
          4472 => x"81",
          4473 => x"17",
          4474 => x"83",
          4475 => x"75",
          4476 => x"f9",
          4477 => x"59",
          4478 => x"08",
          4479 => x"81",
          4480 => x"82",
          4481 => x"59",
          4482 => x"08",
          4483 => x"81",
          4484 => x"07",
          4485 => x"7c",
          4486 => x"ec",
          4487 => x"51",
          4488 => x"81",
          4489 => x"85",
          4490 => x"2e",
          4491 => x"17",
          4492 => x"74",
          4493 => x"73",
          4494 => x"27",
          4495 => x"58",
          4496 => x"80",
          4497 => x"56",
          4498 => x"98",
          4499 => x"26",
          4500 => x"56",
          4501 => x"81",
          4502 => x"52",
          4503 => x"c4",
          4504 => x"ec",
          4505 => x"ba",
          4506 => x"82",
          4507 => x"81",
          4508 => x"06",
          4509 => x"85",
          4510 => x"82",
          4511 => x"09",
          4512 => x"05",
          4513 => x"80",
          4514 => x"07",
          4515 => x"55",
          4516 => x"38",
          4517 => x"09",
          4518 => x"ac",
          4519 => x"80",
          4520 => x"53",
          4521 => x"51",
          4522 => x"82",
          4523 => x"82",
          4524 => x"09",
          4525 => x"82",
          4526 => x"07",
          4527 => x"55",
          4528 => x"2e",
          4529 => x"80",
          4530 => x"75",
          4531 => x"76",
          4532 => x"3f",
          4533 => x"08",
          4534 => x"38",
          4535 => x"0c",
          4536 => x"fe",
          4537 => x"08",
          4538 => x"74",
          4539 => x"ff",
          4540 => x"0c",
          4541 => x"81",
          4542 => x"84",
          4543 => x"39",
          4544 => x"81",
          4545 => x"8c",
          4546 => x"8c",
          4547 => x"ec",
          4548 => x"39",
          4549 => x"55",
          4550 => x"ec",
          4551 => x"0d",
          4552 => x"0d",
          4553 => x"55",
          4554 => x"82",
          4555 => x"58",
          4556 => x"85",
          4557 => x"da",
          4558 => x"74",
          4559 => x"3f",
          4560 => x"08",
          4561 => x"08",
          4562 => x"59",
          4563 => x"77",
          4564 => x"70",
          4565 => x"bb",
          4566 => x"84",
          4567 => x"56",
          4568 => x"58",
          4569 => x"97",
          4570 => x"75",
          4571 => x"52",
          4572 => x"51",
          4573 => x"82",
          4574 => x"80",
          4575 => x"8a",
          4576 => x"32",
          4577 => x"05",
          4578 => x"70",
          4579 => x"51",
          4580 => x"82",
          4581 => x"8a",
          4582 => x"f8",
          4583 => x"7c",
          4584 => x"56",
          4585 => x"80",
          4586 => x"f1",
          4587 => x"06",
          4588 => x"e9",
          4589 => x"18",
          4590 => x"08",
          4591 => x"38",
          4592 => x"82",
          4593 => x"38",
          4594 => x"54",
          4595 => x"74",
          4596 => x"82",
          4597 => x"22",
          4598 => x"79",
          4599 => x"38",
          4600 => x"98",
          4601 => x"cd",
          4602 => x"22",
          4603 => x"54",
          4604 => x"26",
          4605 => x"52",
          4606 => x"a8",
          4607 => x"ec",
          4608 => x"85",
          4609 => x"2e",
          4610 => x"0b",
          4611 => x"08",
          4612 => x"98",
          4613 => x"85",
          4614 => x"85",
          4615 => x"bd",
          4616 => x"31",
          4617 => x"73",
          4618 => x"f4",
          4619 => x"85",
          4620 => x"18",
          4621 => x"18",
          4622 => x"08",
          4623 => x"72",
          4624 => x"38",
          4625 => x"58",
          4626 => x"89",
          4627 => x"18",
          4628 => x"ff",
          4629 => x"05",
          4630 => x"80",
          4631 => x"85",
          4632 => x"3d",
          4633 => x"3d",
          4634 => x"08",
          4635 => x"a0",
          4636 => x"54",
          4637 => x"77",
          4638 => x"80",
          4639 => x"0c",
          4640 => x"53",
          4641 => x"80",
          4642 => x"38",
          4643 => x"06",
          4644 => x"b5",
          4645 => x"98",
          4646 => x"14",
          4647 => x"92",
          4648 => x"2a",
          4649 => x"56",
          4650 => x"26",
          4651 => x"80",
          4652 => x"16",
          4653 => x"77",
          4654 => x"53",
          4655 => x"38",
          4656 => x"51",
          4657 => x"82",
          4658 => x"53",
          4659 => x"0b",
          4660 => x"08",
          4661 => x"38",
          4662 => x"85",
          4663 => x"2e",
          4664 => x"98",
          4665 => x"85",
          4666 => x"80",
          4667 => x"8a",
          4668 => x"15",
          4669 => x"80",
          4670 => x"14",
          4671 => x"51",
          4672 => x"82",
          4673 => x"53",
          4674 => x"85",
          4675 => x"2e",
          4676 => x"82",
          4677 => x"ec",
          4678 => x"ba",
          4679 => x"82",
          4680 => x"ff",
          4681 => x"82",
          4682 => x"52",
          4683 => x"f1",
          4684 => x"ec",
          4685 => x"72",
          4686 => x"72",
          4687 => x"f2",
          4688 => x"85",
          4689 => x"15",
          4690 => x"15",
          4691 => x"b4",
          4692 => x"0c",
          4693 => x"82",
          4694 => x"8a",
          4695 => x"f7",
          4696 => x"7d",
          4697 => x"5b",
          4698 => x"76",
          4699 => x"3f",
          4700 => x"08",
          4701 => x"ec",
          4702 => x"38",
          4703 => x"08",
          4704 => x"08",
          4705 => x"ef",
          4706 => x"85",
          4707 => x"82",
          4708 => x"80",
          4709 => x"85",
          4710 => x"18",
          4711 => x"51",
          4712 => x"81",
          4713 => x"81",
          4714 => x"81",
          4715 => x"ec",
          4716 => x"83",
          4717 => x"77",
          4718 => x"72",
          4719 => x"38",
          4720 => x"75",
          4721 => x"81",
          4722 => x"a5",
          4723 => x"ec",
          4724 => x"52",
          4725 => x"8e",
          4726 => x"ec",
          4727 => x"85",
          4728 => x"2e",
          4729 => x"73",
          4730 => x"81",
          4731 => x"87",
          4732 => x"85",
          4733 => x"3d",
          4734 => x"3d",
          4735 => x"11",
          4736 => x"dd",
          4737 => x"ec",
          4738 => x"ff",
          4739 => x"33",
          4740 => x"71",
          4741 => x"81",
          4742 => x"94",
          4743 => x"c1",
          4744 => x"ec",
          4745 => x"73",
          4746 => x"82",
          4747 => x"85",
          4748 => x"fc",
          4749 => x"79",
          4750 => x"ff",
          4751 => x"12",
          4752 => x"eb",
          4753 => x"70",
          4754 => x"72",
          4755 => x"81",
          4756 => x"73",
          4757 => x"94",
          4758 => x"c7",
          4759 => x"0d",
          4760 => x"0d",
          4761 => x"55",
          4762 => x"5a",
          4763 => x"08",
          4764 => x"8a",
          4765 => x"08",
          4766 => x"ee",
          4767 => x"85",
          4768 => x"82",
          4769 => x"80",
          4770 => x"15",
          4771 => x"55",
          4772 => x"38",
          4773 => x"e6",
          4774 => x"33",
          4775 => x"70",
          4776 => x"58",
          4777 => x"86",
          4778 => x"85",
          4779 => x"73",
          4780 => x"83",
          4781 => x"73",
          4782 => x"38",
          4783 => x"06",
          4784 => x"80",
          4785 => x"75",
          4786 => x"38",
          4787 => x"08",
          4788 => x"54",
          4789 => x"2e",
          4790 => x"83",
          4791 => x"73",
          4792 => x"38",
          4793 => x"51",
          4794 => x"82",
          4795 => x"58",
          4796 => x"08",
          4797 => x"15",
          4798 => x"38",
          4799 => x"0b",
          4800 => x"77",
          4801 => x"0c",
          4802 => x"04",
          4803 => x"77",
          4804 => x"54",
          4805 => x"51",
          4806 => x"82",
          4807 => x"55",
          4808 => x"08",
          4809 => x"14",
          4810 => x"51",
          4811 => x"82",
          4812 => x"55",
          4813 => x"08",
          4814 => x"53",
          4815 => x"08",
          4816 => x"08",
          4817 => x"3f",
          4818 => x"14",
          4819 => x"08",
          4820 => x"3f",
          4821 => x"17",
          4822 => x"85",
          4823 => x"3d",
          4824 => x"3d",
          4825 => x"08",
          4826 => x"54",
          4827 => x"53",
          4828 => x"82",
          4829 => x"8d",
          4830 => x"08",
          4831 => x"34",
          4832 => x"15",
          4833 => x"0d",
          4834 => x"0d",
          4835 => x"57",
          4836 => x"17",
          4837 => x"08",
          4838 => x"82",
          4839 => x"89",
          4840 => x"55",
          4841 => x"14",
          4842 => x"16",
          4843 => x"71",
          4844 => x"38",
          4845 => x"09",
          4846 => x"38",
          4847 => x"73",
          4848 => x"81",
          4849 => x"ae",
          4850 => x"05",
          4851 => x"15",
          4852 => x"70",
          4853 => x"34",
          4854 => x"8a",
          4855 => x"38",
          4856 => x"05",
          4857 => x"81",
          4858 => x"17",
          4859 => x"12",
          4860 => x"34",
          4861 => x"9c",
          4862 => x"e7",
          4863 => x"85",
          4864 => x"0c",
          4865 => x"e7",
          4866 => x"85",
          4867 => x"17",
          4868 => x"51",
          4869 => x"82",
          4870 => x"84",
          4871 => x"3d",
          4872 => x"3d",
          4873 => x"08",
          4874 => x"61",
          4875 => x"55",
          4876 => x"2e",
          4877 => x"55",
          4878 => x"2e",
          4879 => x"80",
          4880 => x"94",
          4881 => x"1c",
          4882 => x"81",
          4883 => x"61",
          4884 => x"56",
          4885 => x"2e",
          4886 => x"83",
          4887 => x"73",
          4888 => x"70",
          4889 => x"70",
          4890 => x"07",
          4891 => x"73",
          4892 => x"88",
          4893 => x"70",
          4894 => x"73",
          4895 => x"38",
          4896 => x"ab",
          4897 => x"52",
          4898 => x"8f",
          4899 => x"ec",
          4900 => x"a6",
          4901 => x"61",
          4902 => x"5a",
          4903 => x"a0",
          4904 => x"e7",
          4905 => x"70",
          4906 => x"79",
          4907 => x"73",
          4908 => x"81",
          4909 => x"38",
          4910 => x"33",
          4911 => x"ae",
          4912 => x"81",
          4913 => x"2a",
          4914 => x"07",
          4915 => x"5a",
          4916 => x"8c",
          4917 => x"54",
          4918 => x"81",
          4919 => x"39",
          4920 => x"70",
          4921 => x"70",
          4922 => x"51",
          4923 => x"dc",
          4924 => x"73",
          4925 => x"38",
          4926 => x"82",
          4927 => x"19",
          4928 => x"54",
          4929 => x"82",
          4930 => x"54",
          4931 => x"78",
          4932 => x"81",
          4933 => x"54",
          4934 => x"82",
          4935 => x"af",
          4936 => x"81",
          4937 => x"dc",
          4938 => x"81",
          4939 => x"25",
          4940 => x"07",
          4941 => x"51",
          4942 => x"2e",
          4943 => x"39",
          4944 => x"80",
          4945 => x"33",
          4946 => x"73",
          4947 => x"81",
          4948 => x"81",
          4949 => x"dc",
          4950 => x"81",
          4951 => x"25",
          4952 => x"51",
          4953 => x"38",
          4954 => x"75",
          4955 => x"81",
          4956 => x"81",
          4957 => x"27",
          4958 => x"73",
          4959 => x"38",
          4960 => x"70",
          4961 => x"77",
          4962 => x"09",
          4963 => x"80",
          4964 => x"2a",
          4965 => x"56",
          4966 => x"81",
          4967 => x"57",
          4968 => x"eb",
          4969 => x"2b",
          4970 => x"25",
          4971 => x"80",
          4972 => x"ff",
          4973 => x"57",
          4974 => x"e6",
          4975 => x"85",
          4976 => x"2e",
          4977 => x"18",
          4978 => x"1a",
          4979 => x"56",
          4980 => x"3f",
          4981 => x"08",
          4982 => x"e8",
          4983 => x"54",
          4984 => x"80",
          4985 => x"17",
          4986 => x"34",
          4987 => x"11",
          4988 => x"74",
          4989 => x"75",
          4990 => x"d4",
          4991 => x"3f",
          4992 => x"08",
          4993 => x"9f",
          4994 => x"99",
          4995 => x"e0",
          4996 => x"ff",
          4997 => x"79",
          4998 => x"74",
          4999 => x"57",
          5000 => x"77",
          5001 => x"76",
          5002 => x"38",
          5003 => x"73",
          5004 => x"09",
          5005 => x"38",
          5006 => x"84",
          5007 => x"27",
          5008 => x"39",
          5009 => x"f2",
          5010 => x"80",
          5011 => x"54",
          5012 => x"34",
          5013 => x"58",
          5014 => x"f2",
          5015 => x"85",
          5016 => x"82",
          5017 => x"80",
          5018 => x"1b",
          5019 => x"51",
          5020 => x"82",
          5021 => x"56",
          5022 => x"08",
          5023 => x"9c",
          5024 => x"33",
          5025 => x"80",
          5026 => x"38",
          5027 => x"bf",
          5028 => x"86",
          5029 => x"15",
          5030 => x"2a",
          5031 => x"51",
          5032 => x"92",
          5033 => x"79",
          5034 => x"e4",
          5035 => x"85",
          5036 => x"2e",
          5037 => x"52",
          5038 => x"aa",
          5039 => x"39",
          5040 => x"33",
          5041 => x"80",
          5042 => x"74",
          5043 => x"81",
          5044 => x"38",
          5045 => x"70",
          5046 => x"82",
          5047 => x"54",
          5048 => x"96",
          5049 => x"06",
          5050 => x"2e",
          5051 => x"ff",
          5052 => x"1c",
          5053 => x"80",
          5054 => x"81",
          5055 => x"ba",
          5056 => x"b6",
          5057 => x"2a",
          5058 => x"51",
          5059 => x"38",
          5060 => x"70",
          5061 => x"81",
          5062 => x"55",
          5063 => x"e1",
          5064 => x"08",
          5065 => x"1d",
          5066 => x"7c",
          5067 => x"3f",
          5068 => x"08",
          5069 => x"fa",
          5070 => x"82",
          5071 => x"8f",
          5072 => x"f6",
          5073 => x"5b",
          5074 => x"70",
          5075 => x"59",
          5076 => x"73",
          5077 => x"cc",
          5078 => x"81",
          5079 => x"70",
          5080 => x"52",
          5081 => x"8d",
          5082 => x"38",
          5083 => x"09",
          5084 => x"ab",
          5085 => x"d0",
          5086 => x"ff",
          5087 => x"53",
          5088 => x"91",
          5089 => x"73",
          5090 => x"d0",
          5091 => x"71",
          5092 => x"fd",
          5093 => x"81",
          5094 => x"55",
          5095 => x"55",
          5096 => x"81",
          5097 => x"74",
          5098 => x"56",
          5099 => x"12",
          5100 => x"70",
          5101 => x"38",
          5102 => x"81",
          5103 => x"51",
          5104 => x"51",
          5105 => x"89",
          5106 => x"70",
          5107 => x"53",
          5108 => x"81",
          5109 => x"2a",
          5110 => x"72",
          5111 => x"06",
          5112 => x"ff",
          5113 => x"09",
          5114 => x"77",
          5115 => x"81",
          5116 => x"07",
          5117 => x"9f",
          5118 => x"54",
          5119 => x"80",
          5120 => x"81",
          5121 => x"59",
          5122 => x"25",
          5123 => x"8b",
          5124 => x"24",
          5125 => x"76",
          5126 => x"78",
          5127 => x"82",
          5128 => x"51",
          5129 => x"ec",
          5130 => x"0d",
          5131 => x"0d",
          5132 => x"0b",
          5133 => x"ff",
          5134 => x"0c",
          5135 => x"51",
          5136 => x"84",
          5137 => x"ec",
          5138 => x"38",
          5139 => x"51",
          5140 => x"82",
          5141 => x"83",
          5142 => x"54",
          5143 => x"82",
          5144 => x"09",
          5145 => x"e5",
          5146 => x"b4",
          5147 => x"57",
          5148 => x"2e",
          5149 => x"83",
          5150 => x"74",
          5151 => x"70",
          5152 => x"70",
          5153 => x"07",
          5154 => x"73",
          5155 => x"81",
          5156 => x"81",
          5157 => x"83",
          5158 => x"e4",
          5159 => x"16",
          5160 => x"3f",
          5161 => x"08",
          5162 => x"ec",
          5163 => x"9d",
          5164 => x"81",
          5165 => x"81",
          5166 => x"df",
          5167 => x"85",
          5168 => x"82",
          5169 => x"80",
          5170 => x"82",
          5171 => x"85",
          5172 => x"3d",
          5173 => x"3d",
          5174 => x"84",
          5175 => x"05",
          5176 => x"80",
          5177 => x"51",
          5178 => x"82",
          5179 => x"58",
          5180 => x"0b",
          5181 => x"08",
          5182 => x"38",
          5183 => x"08",
          5184 => x"9d",
          5185 => x"55",
          5186 => x"73",
          5187 => x"ee",
          5188 => x"0c",
          5189 => x"06",
          5190 => x"57",
          5191 => x"ae",
          5192 => x"33",
          5193 => x"3f",
          5194 => x"08",
          5195 => x"70",
          5196 => x"55",
          5197 => x"76",
          5198 => x"c0",
          5199 => x"2a",
          5200 => x"51",
          5201 => x"72",
          5202 => x"86",
          5203 => x"74",
          5204 => x"15",
          5205 => x"81",
          5206 => x"d7",
          5207 => x"85",
          5208 => x"ff",
          5209 => x"06",
          5210 => x"56",
          5211 => x"38",
          5212 => x"8f",
          5213 => x"2a",
          5214 => x"51",
          5215 => x"72",
          5216 => x"80",
          5217 => x"52",
          5218 => x"3f",
          5219 => x"08",
          5220 => x"57",
          5221 => x"09",
          5222 => x"e2",
          5223 => x"74",
          5224 => x"56",
          5225 => x"33",
          5226 => x"72",
          5227 => x"38",
          5228 => x"51",
          5229 => x"82",
          5230 => x"57",
          5231 => x"84",
          5232 => x"ff",
          5233 => x"56",
          5234 => x"25",
          5235 => x"0b",
          5236 => x"56",
          5237 => x"05",
          5238 => x"83",
          5239 => x"2e",
          5240 => x"52",
          5241 => x"c5",
          5242 => x"ec",
          5243 => x"06",
          5244 => x"27",
          5245 => x"16",
          5246 => x"27",
          5247 => x"56",
          5248 => x"84",
          5249 => x"56",
          5250 => x"84",
          5251 => x"14",
          5252 => x"3f",
          5253 => x"08",
          5254 => x"06",
          5255 => x"80",
          5256 => x"06",
          5257 => x"80",
          5258 => x"db",
          5259 => x"85",
          5260 => x"ff",
          5261 => x"77",
          5262 => x"d8",
          5263 => x"b8",
          5264 => x"ec",
          5265 => x"9c",
          5266 => x"c4",
          5267 => x"15",
          5268 => x"14",
          5269 => x"70",
          5270 => x"51",
          5271 => x"56",
          5272 => x"84",
          5273 => x"81",
          5274 => x"77",
          5275 => x"9a",
          5276 => x"ec",
          5277 => x"15",
          5278 => x"72",
          5279 => x"72",
          5280 => x"38",
          5281 => x"06",
          5282 => x"2e",
          5283 => x"56",
          5284 => x"80",
          5285 => x"da",
          5286 => x"85",
          5287 => x"82",
          5288 => x"88",
          5289 => x"8f",
          5290 => x"56",
          5291 => x"38",
          5292 => x"51",
          5293 => x"82",
          5294 => x"83",
          5295 => x"55",
          5296 => x"80",
          5297 => x"da",
          5298 => x"85",
          5299 => x"80",
          5300 => x"da",
          5301 => x"85",
          5302 => x"ff",
          5303 => x"8d",
          5304 => x"2e",
          5305 => x"88",
          5306 => x"1b",
          5307 => x"05",
          5308 => x"75",
          5309 => x"38",
          5310 => x"52",
          5311 => x"51",
          5312 => x"3f",
          5313 => x"08",
          5314 => x"ec",
          5315 => x"82",
          5316 => x"85",
          5317 => x"ff",
          5318 => x"26",
          5319 => x"57",
          5320 => x"f5",
          5321 => x"82",
          5322 => x"f5",
          5323 => x"81",
          5324 => x"8d",
          5325 => x"2e",
          5326 => x"82",
          5327 => x"16",
          5328 => x"16",
          5329 => x"70",
          5330 => x"7a",
          5331 => x"0c",
          5332 => x"83",
          5333 => x"06",
          5334 => x"de",
          5335 => x"81",
          5336 => x"ec",
          5337 => x"ff",
          5338 => x"56",
          5339 => x"38",
          5340 => x"38",
          5341 => x"51",
          5342 => x"82",
          5343 => x"a8",
          5344 => x"82",
          5345 => x"39",
          5346 => x"80",
          5347 => x"38",
          5348 => x"15",
          5349 => x"53",
          5350 => x"8e",
          5351 => x"75",
          5352 => x"76",
          5353 => x"51",
          5354 => x"ff",
          5355 => x"53",
          5356 => x"9c",
          5357 => x"81",
          5358 => x"0b",
          5359 => x"ff",
          5360 => x"0c",
          5361 => x"84",
          5362 => x"83",
          5363 => x"06",
          5364 => x"80",
          5365 => x"d8",
          5366 => x"85",
          5367 => x"ff",
          5368 => x"72",
          5369 => x"81",
          5370 => x"38",
          5371 => x"73",
          5372 => x"3f",
          5373 => x"08",
          5374 => x"82",
          5375 => x"84",
          5376 => x"b2",
          5377 => x"d9",
          5378 => x"ec",
          5379 => x"ff",
          5380 => x"82",
          5381 => x"09",
          5382 => x"c8",
          5383 => x"51",
          5384 => x"82",
          5385 => x"84",
          5386 => x"d2",
          5387 => x"06",
          5388 => x"98",
          5389 => x"c0",
          5390 => x"ec",
          5391 => x"85",
          5392 => x"09",
          5393 => x"38",
          5394 => x"51",
          5395 => x"82",
          5396 => x"90",
          5397 => x"a0",
          5398 => x"9c",
          5399 => x"ec",
          5400 => x"0c",
          5401 => x"82",
          5402 => x"81",
          5403 => x"82",
          5404 => x"72",
          5405 => x"80",
          5406 => x"0c",
          5407 => x"82",
          5408 => x"91",
          5409 => x"fb",
          5410 => x"54",
          5411 => x"80",
          5412 => x"73",
          5413 => x"80",
          5414 => x"72",
          5415 => x"80",
          5416 => x"86",
          5417 => x"15",
          5418 => x"71",
          5419 => x"81",
          5420 => x"81",
          5421 => x"d0",
          5422 => x"85",
          5423 => x"06",
          5424 => x"38",
          5425 => x"54",
          5426 => x"80",
          5427 => x"71",
          5428 => x"82",
          5429 => x"87",
          5430 => x"fa",
          5431 => x"ab",
          5432 => x"58",
          5433 => x"05",
          5434 => x"d7",
          5435 => x"80",
          5436 => x"ec",
          5437 => x"38",
          5438 => x"08",
          5439 => x"9d",
          5440 => x"08",
          5441 => x"80",
          5442 => x"80",
          5443 => x"54",
          5444 => x"84",
          5445 => x"34",
          5446 => x"75",
          5447 => x"2e",
          5448 => x"53",
          5449 => x"53",
          5450 => x"f7",
          5451 => x"85",
          5452 => x"73",
          5453 => x"0c",
          5454 => x"04",
          5455 => x"67",
          5456 => x"80",
          5457 => x"59",
          5458 => x"78",
          5459 => x"ca",
          5460 => x"06",
          5461 => x"3d",
          5462 => x"99",
          5463 => x"52",
          5464 => x"3f",
          5465 => x"08",
          5466 => x"ec",
          5467 => x"38",
          5468 => x"52",
          5469 => x"52",
          5470 => x"3f",
          5471 => x"08",
          5472 => x"ec",
          5473 => x"02",
          5474 => x"33",
          5475 => x"55",
          5476 => x"25",
          5477 => x"55",
          5478 => x"54",
          5479 => x"81",
          5480 => x"80",
          5481 => x"74",
          5482 => x"81",
          5483 => x"75",
          5484 => x"3f",
          5485 => x"08",
          5486 => x"02",
          5487 => x"91",
          5488 => x"81",
          5489 => x"82",
          5490 => x"06",
          5491 => x"80",
          5492 => x"88",
          5493 => x"39",
          5494 => x"58",
          5495 => x"38",
          5496 => x"70",
          5497 => x"54",
          5498 => x"81",
          5499 => x"52",
          5500 => x"86",
          5501 => x"ec",
          5502 => x"88",
          5503 => x"62",
          5504 => x"d4",
          5505 => x"54",
          5506 => x"15",
          5507 => x"62",
          5508 => x"e8",
          5509 => x"52",
          5510 => x"51",
          5511 => x"7a",
          5512 => x"83",
          5513 => x"80",
          5514 => x"38",
          5515 => x"08",
          5516 => x"53",
          5517 => x"3d",
          5518 => x"dd",
          5519 => x"85",
          5520 => x"82",
          5521 => x"82",
          5522 => x"39",
          5523 => x"38",
          5524 => x"33",
          5525 => x"70",
          5526 => x"55",
          5527 => x"2e",
          5528 => x"55",
          5529 => x"77",
          5530 => x"81",
          5531 => x"73",
          5532 => x"38",
          5533 => x"54",
          5534 => x"a0",
          5535 => x"82",
          5536 => x"52",
          5537 => x"f5",
          5538 => x"ec",
          5539 => x"18",
          5540 => x"55",
          5541 => x"ec",
          5542 => x"38",
          5543 => x"70",
          5544 => x"54",
          5545 => x"86",
          5546 => x"c0",
          5547 => x"b0",
          5548 => x"1b",
          5549 => x"1b",
          5550 => x"70",
          5551 => x"ba",
          5552 => x"ec",
          5553 => x"ec",
          5554 => x"0c",
          5555 => x"52",
          5556 => x"3f",
          5557 => x"08",
          5558 => x"08",
          5559 => x"77",
          5560 => x"86",
          5561 => x"1a",
          5562 => x"1a",
          5563 => x"91",
          5564 => x"0b",
          5565 => x"80",
          5566 => x"0c",
          5567 => x"70",
          5568 => x"54",
          5569 => x"81",
          5570 => x"85",
          5571 => x"2e",
          5572 => x"82",
          5573 => x"94",
          5574 => x"17",
          5575 => x"2b",
          5576 => x"57",
          5577 => x"52",
          5578 => x"f8",
          5579 => x"ec",
          5580 => x"85",
          5581 => x"26",
          5582 => x"55",
          5583 => x"08",
          5584 => x"81",
          5585 => x"79",
          5586 => x"31",
          5587 => x"81",
          5588 => x"07",
          5589 => x"54",
          5590 => x"8a",
          5591 => x"75",
          5592 => x"73",
          5593 => x"98",
          5594 => x"a9",
          5595 => x"ff",
          5596 => x"80",
          5597 => x"76",
          5598 => x"d5",
          5599 => x"85",
          5600 => x"38",
          5601 => x"39",
          5602 => x"82",
          5603 => x"05",
          5604 => x"84",
          5605 => x"0c",
          5606 => x"82",
          5607 => x"97",
          5608 => x"f2",
          5609 => x"63",
          5610 => x"40",
          5611 => x"7e",
          5612 => x"fc",
          5613 => x"51",
          5614 => x"82",
          5615 => x"55",
          5616 => x"08",
          5617 => x"19",
          5618 => x"80",
          5619 => x"74",
          5620 => x"39",
          5621 => x"81",
          5622 => x"56",
          5623 => x"82",
          5624 => x"39",
          5625 => x"1a",
          5626 => x"82",
          5627 => x"0b",
          5628 => x"81",
          5629 => x"39",
          5630 => x"94",
          5631 => x"55",
          5632 => x"83",
          5633 => x"7b",
          5634 => x"89",
          5635 => x"08",
          5636 => x"06",
          5637 => x"81",
          5638 => x"8a",
          5639 => x"05",
          5640 => x"06",
          5641 => x"a8",
          5642 => x"38",
          5643 => x"55",
          5644 => x"19",
          5645 => x"51",
          5646 => x"82",
          5647 => x"55",
          5648 => x"ff",
          5649 => x"ff",
          5650 => x"38",
          5651 => x"0c",
          5652 => x"52",
          5653 => x"9b",
          5654 => x"ec",
          5655 => x"ff",
          5656 => x"85",
          5657 => x"7c",
          5658 => x"57",
          5659 => x"80",
          5660 => x"1a",
          5661 => x"22",
          5662 => x"75",
          5663 => x"38",
          5664 => x"58",
          5665 => x"53",
          5666 => x"1b",
          5667 => x"d8",
          5668 => x"ec",
          5669 => x"38",
          5670 => x"33",
          5671 => x"80",
          5672 => x"b0",
          5673 => x"31",
          5674 => x"27",
          5675 => x"80",
          5676 => x"52",
          5677 => x"77",
          5678 => x"7d",
          5679 => x"b0",
          5680 => x"2b",
          5681 => x"76",
          5682 => x"94",
          5683 => x"ff",
          5684 => x"71",
          5685 => x"7b",
          5686 => x"38",
          5687 => x"19",
          5688 => x"51",
          5689 => x"82",
          5690 => x"fe",
          5691 => x"53",
          5692 => x"83",
          5693 => x"b4",
          5694 => x"51",
          5695 => x"7b",
          5696 => x"08",
          5697 => x"76",
          5698 => x"08",
          5699 => x"0c",
          5700 => x"f3",
          5701 => x"75",
          5702 => x"0c",
          5703 => x"04",
          5704 => x"60",
          5705 => x"40",
          5706 => x"80",
          5707 => x"3d",
          5708 => x"77",
          5709 => x"3f",
          5710 => x"08",
          5711 => x"ec",
          5712 => x"91",
          5713 => x"74",
          5714 => x"38",
          5715 => x"b8",
          5716 => x"33",
          5717 => x"70",
          5718 => x"56",
          5719 => x"74",
          5720 => x"a4",
          5721 => x"82",
          5722 => x"34",
          5723 => x"98",
          5724 => x"91",
          5725 => x"56",
          5726 => x"94",
          5727 => x"11",
          5728 => x"76",
          5729 => x"75",
          5730 => x"80",
          5731 => x"38",
          5732 => x"70",
          5733 => x"56",
          5734 => x"fd",
          5735 => x"11",
          5736 => x"77",
          5737 => x"5c",
          5738 => x"38",
          5739 => x"88",
          5740 => x"74",
          5741 => x"52",
          5742 => x"18",
          5743 => x"51",
          5744 => x"82",
          5745 => x"55",
          5746 => x"08",
          5747 => x"ab",
          5748 => x"2e",
          5749 => x"74",
          5750 => x"95",
          5751 => x"19",
          5752 => x"08",
          5753 => x"88",
          5754 => x"55",
          5755 => x"9c",
          5756 => x"09",
          5757 => x"38",
          5758 => x"91",
          5759 => x"ec",
          5760 => x"38",
          5761 => x"52",
          5762 => x"e7",
          5763 => x"ec",
          5764 => x"fe",
          5765 => x"85",
          5766 => x"7c",
          5767 => x"57",
          5768 => x"80",
          5769 => x"1b",
          5770 => x"22",
          5771 => x"75",
          5772 => x"38",
          5773 => x"59",
          5774 => x"53",
          5775 => x"1a",
          5776 => x"8e",
          5777 => x"ec",
          5778 => x"38",
          5779 => x"08",
          5780 => x"56",
          5781 => x"9b",
          5782 => x"53",
          5783 => x"77",
          5784 => x"7d",
          5785 => x"16",
          5786 => x"3f",
          5787 => x"0b",
          5788 => x"78",
          5789 => x"80",
          5790 => x"18",
          5791 => x"08",
          5792 => x"7e",
          5793 => x"3f",
          5794 => x"08",
          5795 => x"7e",
          5796 => x"0c",
          5797 => x"19",
          5798 => x"08",
          5799 => x"84",
          5800 => x"57",
          5801 => x"27",
          5802 => x"56",
          5803 => x"52",
          5804 => x"c9",
          5805 => x"ec",
          5806 => x"38",
          5807 => x"52",
          5808 => x"83",
          5809 => x"b4",
          5810 => x"a4",
          5811 => x"81",
          5812 => x"34",
          5813 => x"7e",
          5814 => x"0c",
          5815 => x"1a",
          5816 => x"94",
          5817 => x"1b",
          5818 => x"5e",
          5819 => x"27",
          5820 => x"55",
          5821 => x"0c",
          5822 => x"90",
          5823 => x"c0",
          5824 => x"90",
          5825 => x"56",
          5826 => x"ec",
          5827 => x"0d",
          5828 => x"0d",
          5829 => x"fc",
          5830 => x"52",
          5831 => x"3f",
          5832 => x"08",
          5833 => x"ec",
          5834 => x"38",
          5835 => x"70",
          5836 => x"81",
          5837 => x"55",
          5838 => x"80",
          5839 => x"16",
          5840 => x"51",
          5841 => x"82",
          5842 => x"57",
          5843 => x"08",
          5844 => x"a4",
          5845 => x"11",
          5846 => x"55",
          5847 => x"16",
          5848 => x"08",
          5849 => x"75",
          5850 => x"c7",
          5851 => x"08",
          5852 => x"51",
          5853 => x"82",
          5854 => x"52",
          5855 => x"c9",
          5856 => x"52",
          5857 => x"c9",
          5858 => x"54",
          5859 => x"15",
          5860 => x"cc",
          5861 => x"85",
          5862 => x"17",
          5863 => x"06",
          5864 => x"90",
          5865 => x"82",
          5866 => x"8a",
          5867 => x"fc",
          5868 => x"70",
          5869 => x"d9",
          5870 => x"ec",
          5871 => x"85",
          5872 => x"38",
          5873 => x"05",
          5874 => x"f1",
          5875 => x"85",
          5876 => x"82",
          5877 => x"87",
          5878 => x"ec",
          5879 => x"72",
          5880 => x"0c",
          5881 => x"04",
          5882 => x"84",
          5883 => x"d3",
          5884 => x"80",
          5885 => x"ec",
          5886 => x"38",
          5887 => x"08",
          5888 => x"34",
          5889 => x"82",
          5890 => x"83",
          5891 => x"ef",
          5892 => x"53",
          5893 => x"05",
          5894 => x"51",
          5895 => x"82",
          5896 => x"55",
          5897 => x"08",
          5898 => x"76",
          5899 => x"93",
          5900 => x"51",
          5901 => x"82",
          5902 => x"55",
          5903 => x"08",
          5904 => x"80",
          5905 => x"70",
          5906 => x"56",
          5907 => x"89",
          5908 => x"94",
          5909 => x"b2",
          5910 => x"05",
          5911 => x"2a",
          5912 => x"51",
          5913 => x"80",
          5914 => x"76",
          5915 => x"52",
          5916 => x"3f",
          5917 => x"08",
          5918 => x"8e",
          5919 => x"ec",
          5920 => x"09",
          5921 => x"38",
          5922 => x"82",
          5923 => x"93",
          5924 => x"e4",
          5925 => x"6f",
          5926 => x"7a",
          5927 => x"9e",
          5928 => x"05",
          5929 => x"51",
          5930 => x"82",
          5931 => x"57",
          5932 => x"08",
          5933 => x"7b",
          5934 => x"94",
          5935 => x"55",
          5936 => x"73",
          5937 => x"ed",
          5938 => x"93",
          5939 => x"55",
          5940 => x"82",
          5941 => x"57",
          5942 => x"08",
          5943 => x"68",
          5944 => x"c9",
          5945 => x"85",
          5946 => x"82",
          5947 => x"82",
          5948 => x"52",
          5949 => x"82",
          5950 => x"ec",
          5951 => x"52",
          5952 => x"97",
          5953 => x"ec",
          5954 => x"85",
          5955 => x"a1",
          5956 => x"74",
          5957 => x"3f",
          5958 => x"08",
          5959 => x"ec",
          5960 => x"69",
          5961 => x"d9",
          5962 => x"82",
          5963 => x"2e",
          5964 => x"52",
          5965 => x"ae",
          5966 => x"ec",
          5967 => x"85",
          5968 => x"2e",
          5969 => x"84",
          5970 => x"06",
          5971 => x"57",
          5972 => x"76",
          5973 => x"9e",
          5974 => x"05",
          5975 => x"dc",
          5976 => x"90",
          5977 => x"81",
          5978 => x"56",
          5979 => x"80",
          5980 => x"02",
          5981 => x"81",
          5982 => x"70",
          5983 => x"56",
          5984 => x"81",
          5985 => x"78",
          5986 => x"38",
          5987 => x"99",
          5988 => x"81",
          5989 => x"18",
          5990 => x"18",
          5991 => x"58",
          5992 => x"33",
          5993 => x"ee",
          5994 => x"6f",
          5995 => x"af",
          5996 => x"8d",
          5997 => x"2e",
          5998 => x"8a",
          5999 => x"6f",
          6000 => x"af",
          6001 => x"0b",
          6002 => x"33",
          6003 => x"81",
          6004 => x"08",
          6005 => x"5c",
          6006 => x"73",
          6007 => x"38",
          6008 => x"1a",
          6009 => x"55",
          6010 => x"38",
          6011 => x"73",
          6012 => x"38",
          6013 => x"76",
          6014 => x"74",
          6015 => x"33",
          6016 => x"05",
          6017 => x"15",
          6018 => x"ba",
          6019 => x"05",
          6020 => x"ff",
          6021 => x"06",
          6022 => x"57",
          6023 => x"18",
          6024 => x"54",
          6025 => x"70",
          6026 => x"34",
          6027 => x"ee",
          6028 => x"34",
          6029 => x"ec",
          6030 => x"0d",
          6031 => x"0d",
          6032 => x"3d",
          6033 => x"71",
          6034 => x"ec",
          6035 => x"85",
          6036 => x"82",
          6037 => x"82",
          6038 => x"15",
          6039 => x"82",
          6040 => x"15",
          6041 => x"76",
          6042 => x"90",
          6043 => x"81",
          6044 => x"06",
          6045 => x"72",
          6046 => x"56",
          6047 => x"54",
          6048 => x"17",
          6049 => x"78",
          6050 => x"38",
          6051 => x"22",
          6052 => x"59",
          6053 => x"78",
          6054 => x"76",
          6055 => x"51",
          6056 => x"3f",
          6057 => x"08",
          6058 => x"54",
          6059 => x"53",
          6060 => x"3f",
          6061 => x"08",
          6062 => x"38",
          6063 => x"05",
          6064 => x"70",
          6065 => x"77",
          6066 => x"18",
          6067 => x"51",
          6068 => x"88",
          6069 => x"73",
          6070 => x"52",
          6071 => x"a0",
          6072 => x"ec",
          6073 => x"85",
          6074 => x"2e",
          6075 => x"82",
          6076 => x"ff",
          6077 => x"38",
          6078 => x"08",
          6079 => x"73",
          6080 => x"73",
          6081 => x"9c",
          6082 => x"27",
          6083 => x"75",
          6084 => x"16",
          6085 => x"17",
          6086 => x"33",
          6087 => x"70",
          6088 => x"55",
          6089 => x"80",
          6090 => x"73",
          6091 => x"cc",
          6092 => x"85",
          6093 => x"82",
          6094 => x"94",
          6095 => x"ec",
          6096 => x"39",
          6097 => x"51",
          6098 => x"82",
          6099 => x"54",
          6100 => x"be",
          6101 => x"27",
          6102 => x"53",
          6103 => x"08",
          6104 => x"73",
          6105 => x"ff",
          6106 => x"15",
          6107 => x"16",
          6108 => x"ff",
          6109 => x"80",
          6110 => x"73",
          6111 => x"c5",
          6112 => x"85",
          6113 => x"38",
          6114 => x"16",
          6115 => x"80",
          6116 => x"0b",
          6117 => x"81",
          6118 => x"75",
          6119 => x"85",
          6120 => x"58",
          6121 => x"54",
          6122 => x"74",
          6123 => x"73",
          6124 => x"90",
          6125 => x"c0",
          6126 => x"90",
          6127 => x"83",
          6128 => x"72",
          6129 => x"38",
          6130 => x"08",
          6131 => x"77",
          6132 => x"80",
          6133 => x"85",
          6134 => x"3d",
          6135 => x"3d",
          6136 => x"89",
          6137 => x"2e",
          6138 => x"80",
          6139 => x"fc",
          6140 => x"3d",
          6141 => x"e1",
          6142 => x"85",
          6143 => x"82",
          6144 => x"80",
          6145 => x"76",
          6146 => x"75",
          6147 => x"3f",
          6148 => x"08",
          6149 => x"ec",
          6150 => x"38",
          6151 => x"70",
          6152 => x"57",
          6153 => x"a2",
          6154 => x"33",
          6155 => x"70",
          6156 => x"55",
          6157 => x"2e",
          6158 => x"16",
          6159 => x"51",
          6160 => x"82",
          6161 => x"88",
          6162 => x"54",
          6163 => x"84",
          6164 => x"52",
          6165 => x"c3",
          6166 => x"ec",
          6167 => x"84",
          6168 => x"06",
          6169 => x"55",
          6170 => x"80",
          6171 => x"80",
          6172 => x"54",
          6173 => x"ec",
          6174 => x"0d",
          6175 => x"0d",
          6176 => x"fc",
          6177 => x"52",
          6178 => x"3f",
          6179 => x"08",
          6180 => x"85",
          6181 => x"0c",
          6182 => x"04",
          6183 => x"77",
          6184 => x"fc",
          6185 => x"53",
          6186 => x"db",
          6187 => x"ec",
          6188 => x"85",
          6189 => x"e1",
          6190 => x"38",
          6191 => x"08",
          6192 => x"cd",
          6193 => x"85",
          6194 => x"80",
          6195 => x"85",
          6196 => x"73",
          6197 => x"3f",
          6198 => x"08",
          6199 => x"ec",
          6200 => x"09",
          6201 => x"38",
          6202 => x"39",
          6203 => x"08",
          6204 => x"52",
          6205 => x"91",
          6206 => x"73",
          6207 => x"3f",
          6208 => x"08",
          6209 => x"09",
          6210 => x"72",
          6211 => x"70",
          6212 => x"08",
          6213 => x"54",
          6214 => x"85",
          6215 => x"3d",
          6216 => x"3d",
          6217 => x"80",
          6218 => x"70",
          6219 => x"52",
          6220 => x"3f",
          6221 => x"08",
          6222 => x"ec",
          6223 => x"64",
          6224 => x"d5",
          6225 => x"85",
          6226 => x"82",
          6227 => x"a0",
          6228 => x"cb",
          6229 => x"98",
          6230 => x"73",
          6231 => x"38",
          6232 => x"39",
          6233 => x"88",
          6234 => x"75",
          6235 => x"3f",
          6236 => x"ec",
          6237 => x"0d",
          6238 => x"0d",
          6239 => x"5c",
          6240 => x"3d",
          6241 => x"93",
          6242 => x"ca",
          6243 => x"ec",
          6244 => x"85",
          6245 => x"87",
          6246 => x"0c",
          6247 => x"11",
          6248 => x"90",
          6249 => x"56",
          6250 => x"74",
          6251 => x"75",
          6252 => x"eb",
          6253 => x"81",
          6254 => x"5b",
          6255 => x"82",
          6256 => x"75",
          6257 => x"73",
          6258 => x"81",
          6259 => x"38",
          6260 => x"57",
          6261 => x"3d",
          6262 => x"c1",
          6263 => x"85",
          6264 => x"2e",
          6265 => x"85",
          6266 => x"2e",
          6267 => x"85",
          6268 => x"81",
          6269 => x"85",
          6270 => x"80",
          6271 => x"81",
          6272 => x"59",
          6273 => x"14",
          6274 => x"c8",
          6275 => x"39",
          6276 => x"82",
          6277 => x"57",
          6278 => x"38",
          6279 => x"18",
          6280 => x"ff",
          6281 => x"82",
          6282 => x"5b",
          6283 => x"08",
          6284 => x"7c",
          6285 => x"12",
          6286 => x"52",
          6287 => x"82",
          6288 => x"06",
          6289 => x"14",
          6290 => x"95",
          6291 => x"ec",
          6292 => x"ff",
          6293 => x"81",
          6294 => x"25",
          6295 => x"59",
          6296 => x"9d",
          6297 => x"51",
          6298 => x"3f",
          6299 => x"08",
          6300 => x"70",
          6301 => x"70",
          6302 => x"84",
          6303 => x"51",
          6304 => x"ff",
          6305 => x"56",
          6306 => x"38",
          6307 => x"7c",
          6308 => x"0c",
          6309 => x"81",
          6310 => x"74",
          6311 => x"7a",
          6312 => x"0c",
          6313 => x"04",
          6314 => x"79",
          6315 => x"05",
          6316 => x"57",
          6317 => x"82",
          6318 => x"56",
          6319 => x"08",
          6320 => x"91",
          6321 => x"75",
          6322 => x"90",
          6323 => x"81",
          6324 => x"06",
          6325 => x"87",
          6326 => x"2e",
          6327 => x"94",
          6328 => x"73",
          6329 => x"27",
          6330 => x"73",
          6331 => x"85",
          6332 => x"88",
          6333 => x"76",
          6334 => x"3f",
          6335 => x"08",
          6336 => x"0c",
          6337 => x"39",
          6338 => x"52",
          6339 => x"bf",
          6340 => x"85",
          6341 => x"2e",
          6342 => x"83",
          6343 => x"82",
          6344 => x"81",
          6345 => x"06",
          6346 => x"56",
          6347 => x"a0",
          6348 => x"82",
          6349 => x"98",
          6350 => x"94",
          6351 => x"08",
          6352 => x"ec",
          6353 => x"51",
          6354 => x"82",
          6355 => x"56",
          6356 => x"8c",
          6357 => x"17",
          6358 => x"07",
          6359 => x"18",
          6360 => x"2e",
          6361 => x"91",
          6362 => x"55",
          6363 => x"ec",
          6364 => x"0d",
          6365 => x"0d",
          6366 => x"3d",
          6367 => x"52",
          6368 => x"da",
          6369 => x"85",
          6370 => x"82",
          6371 => x"81",
          6372 => x"45",
          6373 => x"52",
          6374 => x"52",
          6375 => x"3f",
          6376 => x"08",
          6377 => x"ec",
          6378 => x"38",
          6379 => x"05",
          6380 => x"2a",
          6381 => x"51",
          6382 => x"55",
          6383 => x"38",
          6384 => x"54",
          6385 => x"81",
          6386 => x"80",
          6387 => x"70",
          6388 => x"54",
          6389 => x"81",
          6390 => x"52",
          6391 => x"9a",
          6392 => x"ec",
          6393 => x"2a",
          6394 => x"51",
          6395 => x"80",
          6396 => x"38",
          6397 => x"85",
          6398 => x"15",
          6399 => x"88",
          6400 => x"82",
          6401 => x"5c",
          6402 => x"3d",
          6403 => x"c7",
          6404 => x"85",
          6405 => x"82",
          6406 => x"80",
          6407 => x"85",
          6408 => x"73",
          6409 => x"3f",
          6410 => x"08",
          6411 => x"ec",
          6412 => x"87",
          6413 => x"39",
          6414 => x"08",
          6415 => x"38",
          6416 => x"08",
          6417 => x"77",
          6418 => x"3f",
          6419 => x"08",
          6420 => x"08",
          6421 => x"70",
          6422 => x"08",
          6423 => x"51",
          6424 => x"80",
          6425 => x"73",
          6426 => x"38",
          6427 => x"52",
          6428 => x"e0",
          6429 => x"ec",
          6430 => x"8c",
          6431 => x"ff",
          6432 => x"82",
          6433 => x"55",
          6434 => x"ec",
          6435 => x"0d",
          6436 => x"0d",
          6437 => x"3d",
          6438 => x"9a",
          6439 => x"b6",
          6440 => x"ec",
          6441 => x"85",
          6442 => x"b0",
          6443 => x"69",
          6444 => x"70",
          6445 => x"ea",
          6446 => x"ec",
          6447 => x"85",
          6448 => x"38",
          6449 => x"94",
          6450 => x"ec",
          6451 => x"09",
          6452 => x"88",
          6453 => x"df",
          6454 => x"85",
          6455 => x"51",
          6456 => x"74",
          6457 => x"78",
          6458 => x"8a",
          6459 => x"57",
          6460 => x"82",
          6461 => x"75",
          6462 => x"85",
          6463 => x"38",
          6464 => x"85",
          6465 => x"2e",
          6466 => x"83",
          6467 => x"82",
          6468 => x"ff",
          6469 => x"06",
          6470 => x"54",
          6471 => x"73",
          6472 => x"82",
          6473 => x"52",
          6474 => x"f5",
          6475 => x"ec",
          6476 => x"85",
          6477 => x"9a",
          6478 => x"a0",
          6479 => x"51",
          6480 => x"3f",
          6481 => x"0b",
          6482 => x"78",
          6483 => x"bf",
          6484 => x"88",
          6485 => x"80",
          6486 => x"ff",
          6487 => x"75",
          6488 => x"11",
          6489 => x"cb",
          6490 => x"78",
          6491 => x"80",
          6492 => x"ff",
          6493 => x"78",
          6494 => x"80",
          6495 => x"7f",
          6496 => x"d4",
          6497 => x"c9",
          6498 => x"54",
          6499 => x"15",
          6500 => x"ca",
          6501 => x"85",
          6502 => x"82",
          6503 => x"b2",
          6504 => x"b2",
          6505 => x"96",
          6506 => x"b5",
          6507 => x"53",
          6508 => x"51",
          6509 => x"64",
          6510 => x"8b",
          6511 => x"54",
          6512 => x"15",
          6513 => x"ff",
          6514 => x"82",
          6515 => x"54",
          6516 => x"53",
          6517 => x"51",
          6518 => x"3f",
          6519 => x"ec",
          6520 => x"0d",
          6521 => x"0d",
          6522 => x"05",
          6523 => x"3f",
          6524 => x"3d",
          6525 => x"52",
          6526 => x"d5",
          6527 => x"85",
          6528 => x"82",
          6529 => x"82",
          6530 => x"4d",
          6531 => x"52",
          6532 => x"52",
          6533 => x"3f",
          6534 => x"08",
          6535 => x"ec",
          6536 => x"38",
          6537 => x"05",
          6538 => x"06",
          6539 => x"73",
          6540 => x"a0",
          6541 => x"08",
          6542 => x"ff",
          6543 => x"ff",
          6544 => x"ac",
          6545 => x"92",
          6546 => x"54",
          6547 => x"3f",
          6548 => x"52",
          6549 => x"ca",
          6550 => x"ec",
          6551 => x"85",
          6552 => x"38",
          6553 => x"09",
          6554 => x"38",
          6555 => x"08",
          6556 => x"88",
          6557 => x"39",
          6558 => x"08",
          6559 => x"81",
          6560 => x"38",
          6561 => x"84",
          6562 => x"ec",
          6563 => x"85",
          6564 => x"c8",
          6565 => x"93",
          6566 => x"ff",
          6567 => x"8d",
          6568 => x"b3",
          6569 => x"af",
          6570 => x"17",
          6571 => x"33",
          6572 => x"70",
          6573 => x"55",
          6574 => x"38",
          6575 => x"54",
          6576 => x"34",
          6577 => x"0b",
          6578 => x"8b",
          6579 => x"84",
          6580 => x"06",
          6581 => x"73",
          6582 => x"e5",
          6583 => x"2e",
          6584 => x"75",
          6585 => x"c6",
          6586 => x"85",
          6587 => x"78",
          6588 => x"ff",
          6589 => x"82",
          6590 => x"80",
          6591 => x"38",
          6592 => x"08",
          6593 => x"ff",
          6594 => x"82",
          6595 => x"79",
          6596 => x"58",
          6597 => x"85",
          6598 => x"c0",
          6599 => x"33",
          6600 => x"2e",
          6601 => x"99",
          6602 => x"75",
          6603 => x"c6",
          6604 => x"54",
          6605 => x"15",
          6606 => x"82",
          6607 => x"9c",
          6608 => x"c8",
          6609 => x"85",
          6610 => x"82",
          6611 => x"8c",
          6612 => x"ff",
          6613 => x"82",
          6614 => x"55",
          6615 => x"ec",
          6616 => x"0d",
          6617 => x"0d",
          6618 => x"05",
          6619 => x"05",
          6620 => x"33",
          6621 => x"53",
          6622 => x"05",
          6623 => x"51",
          6624 => x"82",
          6625 => x"55",
          6626 => x"08",
          6627 => x"78",
          6628 => x"95",
          6629 => x"51",
          6630 => x"82",
          6631 => x"55",
          6632 => x"08",
          6633 => x"80",
          6634 => x"81",
          6635 => x"86",
          6636 => x"38",
          6637 => x"61",
          6638 => x"12",
          6639 => x"7a",
          6640 => x"51",
          6641 => x"74",
          6642 => x"78",
          6643 => x"83",
          6644 => x"51",
          6645 => x"3f",
          6646 => x"08",
          6647 => x"85",
          6648 => x"3d",
          6649 => x"3d",
          6650 => x"82",
          6651 => x"d0",
          6652 => x"3d",
          6653 => x"3f",
          6654 => x"08",
          6655 => x"ec",
          6656 => x"38",
          6657 => x"52",
          6658 => x"05",
          6659 => x"3f",
          6660 => x"08",
          6661 => x"ec",
          6662 => x"02",
          6663 => x"33",
          6664 => x"54",
          6665 => x"a6",
          6666 => x"22",
          6667 => x"71",
          6668 => x"53",
          6669 => x"51",
          6670 => x"3f",
          6671 => x"0b",
          6672 => x"76",
          6673 => x"fc",
          6674 => x"ec",
          6675 => x"82",
          6676 => x"93",
          6677 => x"ea",
          6678 => x"6b",
          6679 => x"53",
          6680 => x"05",
          6681 => x"51",
          6682 => x"82",
          6683 => x"82",
          6684 => x"09",
          6685 => x"82",
          6686 => x"07",
          6687 => x"55",
          6688 => x"2e",
          6689 => x"81",
          6690 => x"55",
          6691 => x"2e",
          6692 => x"7b",
          6693 => x"80",
          6694 => x"70",
          6695 => x"bd",
          6696 => x"85",
          6697 => x"82",
          6698 => x"80",
          6699 => x"52",
          6700 => x"ad",
          6701 => x"ec",
          6702 => x"85",
          6703 => x"38",
          6704 => x"08",
          6705 => x"08",
          6706 => x"56",
          6707 => x"19",
          6708 => x"59",
          6709 => x"74",
          6710 => x"56",
          6711 => x"ec",
          6712 => x"75",
          6713 => x"74",
          6714 => x"2e",
          6715 => x"16",
          6716 => x"33",
          6717 => x"73",
          6718 => x"38",
          6719 => x"84",
          6720 => x"06",
          6721 => x"7a",
          6722 => x"76",
          6723 => x"70",
          6724 => x"25",
          6725 => x"80",
          6726 => x"38",
          6727 => x"bc",
          6728 => x"11",
          6729 => x"ff",
          6730 => x"82",
          6731 => x"57",
          6732 => x"08",
          6733 => x"70",
          6734 => x"80",
          6735 => x"83",
          6736 => x"80",
          6737 => x"84",
          6738 => x"a7",
          6739 => x"b4",
          6740 => x"ad",
          6741 => x"85",
          6742 => x"0c",
          6743 => x"ec",
          6744 => x"0d",
          6745 => x"0d",
          6746 => x"3d",
          6747 => x"52",
          6748 => x"ce",
          6749 => x"85",
          6750 => x"85",
          6751 => x"54",
          6752 => x"08",
          6753 => x"8b",
          6754 => x"8b",
          6755 => x"59",
          6756 => x"3f",
          6757 => x"33",
          6758 => x"06",
          6759 => x"57",
          6760 => x"81",
          6761 => x"58",
          6762 => x"06",
          6763 => x"4e",
          6764 => x"ff",
          6765 => x"82",
          6766 => x"80",
          6767 => x"6c",
          6768 => x"53",
          6769 => x"ae",
          6770 => x"85",
          6771 => x"2e",
          6772 => x"88",
          6773 => x"6d",
          6774 => x"55",
          6775 => x"85",
          6776 => x"ff",
          6777 => x"83",
          6778 => x"51",
          6779 => x"26",
          6780 => x"15",
          6781 => x"ff",
          6782 => x"80",
          6783 => x"87",
          6784 => x"b4",
          6785 => x"74",
          6786 => x"38",
          6787 => x"80",
          6788 => x"ad",
          6789 => x"85",
          6790 => x"38",
          6791 => x"27",
          6792 => x"89",
          6793 => x"8b",
          6794 => x"27",
          6795 => x"55",
          6796 => x"81",
          6797 => x"8f",
          6798 => x"2a",
          6799 => x"70",
          6800 => x"34",
          6801 => x"74",
          6802 => x"05",
          6803 => x"17",
          6804 => x"70",
          6805 => x"52",
          6806 => x"73",
          6807 => x"c8",
          6808 => x"33",
          6809 => x"73",
          6810 => x"81",
          6811 => x"80",
          6812 => x"02",
          6813 => x"76",
          6814 => x"51",
          6815 => x"2e",
          6816 => x"87",
          6817 => x"57",
          6818 => x"79",
          6819 => x"80",
          6820 => x"70",
          6821 => x"ba",
          6822 => x"85",
          6823 => x"82",
          6824 => x"80",
          6825 => x"52",
          6826 => x"bf",
          6827 => x"85",
          6828 => x"82",
          6829 => x"8d",
          6830 => x"c4",
          6831 => x"e5",
          6832 => x"c6",
          6833 => x"ec",
          6834 => x"09",
          6835 => x"cc",
          6836 => x"76",
          6837 => x"c4",
          6838 => x"74",
          6839 => x"ff",
          6840 => x"ec",
          6841 => x"85",
          6842 => x"38",
          6843 => x"85",
          6844 => x"67",
          6845 => x"9b",
          6846 => x"88",
          6847 => x"34",
          6848 => x"52",
          6849 => x"aa",
          6850 => x"54",
          6851 => x"15",
          6852 => x"ff",
          6853 => x"82",
          6854 => x"54",
          6855 => x"82",
          6856 => x"9c",
          6857 => x"f2",
          6858 => x"62",
          6859 => x"80",
          6860 => x"93",
          6861 => x"55",
          6862 => x"5e",
          6863 => x"3f",
          6864 => x"08",
          6865 => x"ec",
          6866 => x"38",
          6867 => x"58",
          6868 => x"38",
          6869 => x"97",
          6870 => x"08",
          6871 => x"38",
          6872 => x"70",
          6873 => x"81",
          6874 => x"55",
          6875 => x"87",
          6876 => x"39",
          6877 => x"92",
          6878 => x"82",
          6879 => x"8a",
          6880 => x"89",
          6881 => x"7f",
          6882 => x"56",
          6883 => x"3f",
          6884 => x"06",
          6885 => x"05",
          6886 => x"9f",
          6887 => x"ec",
          6888 => x"19",
          6889 => x"5a",
          6890 => x"81",
          6891 => x"38",
          6892 => x"77",
          6893 => x"82",
          6894 => x"56",
          6895 => x"74",
          6896 => x"ff",
          6897 => x"81",
          6898 => x"55",
          6899 => x"75",
          6900 => x"82",
          6901 => x"ec",
          6902 => x"ff",
          6903 => x"85",
          6904 => x"2e",
          6905 => x"82",
          6906 => x"8e",
          6907 => x"56",
          6908 => x"09",
          6909 => x"38",
          6910 => x"59",
          6911 => x"77",
          6912 => x"06",
          6913 => x"87",
          6914 => x"39",
          6915 => x"ba",
          6916 => x"55",
          6917 => x"2e",
          6918 => x"15",
          6919 => x"2e",
          6920 => x"83",
          6921 => x"75",
          6922 => x"7e",
          6923 => x"ed",
          6924 => x"ec",
          6925 => x"85",
          6926 => x"ce",
          6927 => x"16",
          6928 => x"56",
          6929 => x"38",
          6930 => x"19",
          6931 => x"8c",
          6932 => x"7d",
          6933 => x"38",
          6934 => x"0c",
          6935 => x"0c",
          6936 => x"80",
          6937 => x"73",
          6938 => x"98",
          6939 => x"05",
          6940 => x"57",
          6941 => x"26",
          6942 => x"7b",
          6943 => x"0c",
          6944 => x"81",
          6945 => x"84",
          6946 => x"54",
          6947 => x"ec",
          6948 => x"0d",
          6949 => x"0d",
          6950 => x"88",
          6951 => x"05",
          6952 => x"54",
          6953 => x"c5",
          6954 => x"56",
          6955 => x"85",
          6956 => x"8c",
          6957 => x"85",
          6958 => x"2b",
          6959 => x"11",
          6960 => x"74",
          6961 => x"38",
          6962 => x"82",
          6963 => x"81",
          6964 => x"81",
          6965 => x"ff",
          6966 => x"82",
          6967 => x"81",
          6968 => x"81",
          6969 => x"83",
          6970 => x"cb",
          6971 => x"2a",
          6972 => x"51",
          6973 => x"74",
          6974 => x"99",
          6975 => x"53",
          6976 => x"51",
          6977 => x"3f",
          6978 => x"08",
          6979 => x"55",
          6980 => x"92",
          6981 => x"80",
          6982 => x"38",
          6983 => x"06",
          6984 => x"2e",
          6985 => x"48",
          6986 => x"87",
          6987 => x"79",
          6988 => x"78",
          6989 => x"26",
          6990 => x"19",
          6991 => x"74",
          6992 => x"38",
          6993 => x"ef",
          6994 => x"2a",
          6995 => x"70",
          6996 => x"59",
          6997 => x"7a",
          6998 => x"56",
          6999 => x"05",
          7000 => x"77",
          7001 => x"91",
          7002 => x"cb",
          7003 => x"f8",
          7004 => x"52",
          7005 => x"a3",
          7006 => x"56",
          7007 => x"08",
          7008 => x"77",
          7009 => x"77",
          7010 => x"ec",
          7011 => x"45",
          7012 => x"bf",
          7013 => x"8e",
          7014 => x"26",
          7015 => x"74",
          7016 => x"48",
          7017 => x"75",
          7018 => x"38",
          7019 => x"81",
          7020 => x"83",
          7021 => x"2a",
          7022 => x"56",
          7023 => x"2e",
          7024 => x"87",
          7025 => x"82",
          7026 => x"38",
          7027 => x"55",
          7028 => x"83",
          7029 => x"81",
          7030 => x"56",
          7031 => x"80",
          7032 => x"38",
          7033 => x"83",
          7034 => x"06",
          7035 => x"78",
          7036 => x"91",
          7037 => x"0b",
          7038 => x"22",
          7039 => x"80",
          7040 => x"74",
          7041 => x"38",
          7042 => x"56",
          7043 => x"17",
          7044 => x"57",
          7045 => x"2e",
          7046 => x"75",
          7047 => x"79",
          7048 => x"fe",
          7049 => x"82",
          7050 => x"82",
          7051 => x"11",
          7052 => x"55",
          7053 => x"0b",
          7054 => x"08",
          7055 => x"05",
          7056 => x"ff",
          7057 => x"27",
          7058 => x"88",
          7059 => x"ae",
          7060 => x"2a",
          7061 => x"82",
          7062 => x"56",
          7063 => x"2e",
          7064 => x"77",
          7065 => x"82",
          7066 => x"79",
          7067 => x"70",
          7068 => x"5a",
          7069 => x"86",
          7070 => x"27",
          7071 => x"52",
          7072 => x"c1",
          7073 => x"85",
          7074 => x"85",
          7075 => x"84",
          7076 => x"85",
          7077 => x"f5",
          7078 => x"81",
          7079 => x"ec",
          7080 => x"82",
          7081 => x"11",
          7082 => x"2a",
          7083 => x"51",
          7084 => x"ff",
          7085 => x"5d",
          7086 => x"44",
          7087 => x"11",
          7088 => x"70",
          7089 => x"71",
          7090 => x"70",
          7091 => x"31",
          7092 => x"57",
          7093 => x"83",
          7094 => x"06",
          7095 => x"1c",
          7096 => x"5c",
          7097 => x"1d",
          7098 => x"2b",
          7099 => x"31",
          7100 => x"55",
          7101 => x"87",
          7102 => x"7c",
          7103 => x"7a",
          7104 => x"31",
          7105 => x"c0",
          7106 => x"85",
          7107 => x"7d",
          7108 => x"81",
          7109 => x"82",
          7110 => x"83",
          7111 => x"80",
          7112 => x"87",
          7113 => x"81",
          7114 => x"fd",
          7115 => x"fa",
          7116 => x"2e",
          7117 => x"80",
          7118 => x"ff",
          7119 => x"85",
          7120 => x"a0",
          7121 => x"38",
          7122 => x"74",
          7123 => x"86",
          7124 => x"fd",
          7125 => x"81",
          7126 => x"80",
          7127 => x"83",
          7128 => x"39",
          7129 => x"08",
          7130 => x"92",
          7131 => x"ba",
          7132 => x"59",
          7133 => x"27",
          7134 => x"86",
          7135 => x"55",
          7136 => x"09",
          7137 => x"38",
          7138 => x"f5",
          7139 => x"38",
          7140 => x"55",
          7141 => x"86",
          7142 => x"80",
          7143 => x"7a",
          7144 => x"ef",
          7145 => x"81",
          7146 => x"7a",
          7147 => x"c0",
          7148 => x"52",
          7149 => x"ff",
          7150 => x"79",
          7151 => x"7b",
          7152 => x"06",
          7153 => x"51",
          7154 => x"3f",
          7155 => x"1c",
          7156 => x"32",
          7157 => x"05",
          7158 => x"84",
          7159 => x"51",
          7160 => x"51",
          7161 => x"3f",
          7162 => x"83",
          7163 => x"90",
          7164 => x"ff",
          7165 => x"93",
          7166 => x"a0",
          7167 => x"39",
          7168 => x"1b",
          7169 => x"b9",
          7170 => x"95",
          7171 => x"52",
          7172 => x"ff",
          7173 => x"81",
          7174 => x"1b",
          7175 => x"83",
          7176 => x"9c",
          7177 => x"a0",
          7178 => x"83",
          7179 => x"06",
          7180 => x"82",
          7181 => x"52",
          7182 => x"51",
          7183 => x"3f",
          7184 => x"1b",
          7185 => x"f9",
          7186 => x"ac",
          7187 => x"9f",
          7188 => x"52",
          7189 => x"ff",
          7190 => x"86",
          7191 => x"51",
          7192 => x"3f",
          7193 => x"80",
          7194 => x"a9",
          7195 => x"1c",
          7196 => x"81",
          7197 => x"80",
          7198 => x"ae",
          7199 => x"b2",
          7200 => x"1b",
          7201 => x"b9",
          7202 => x"ff",
          7203 => x"96",
          7204 => x"9f",
          7205 => x"80",
          7206 => x"34",
          7207 => x"1c",
          7208 => x"81",
          7209 => x"ab",
          7210 => x"9f",
          7211 => x"d4",
          7212 => x"fe",
          7213 => x"59",
          7214 => x"3f",
          7215 => x"53",
          7216 => x"51",
          7217 => x"3f",
          7218 => x"85",
          7219 => x"e7",
          7220 => x"2e",
          7221 => x"80",
          7222 => x"54",
          7223 => x"53",
          7224 => x"51",
          7225 => x"3f",
          7226 => x"80",
          7227 => x"ff",
          7228 => x"84",
          7229 => x"d2",
          7230 => x"ff",
          7231 => x"86",
          7232 => x"f2",
          7233 => x"1b",
          7234 => x"b5",
          7235 => x"52",
          7236 => x"51",
          7237 => x"3f",
          7238 => x"ec",
          7239 => x"9e",
          7240 => x"d4",
          7241 => x"51",
          7242 => x"3f",
          7243 => x"87",
          7244 => x"52",
          7245 => x"9a",
          7246 => x"54",
          7247 => x"7a",
          7248 => x"ff",
          7249 => x"65",
          7250 => x"7a",
          7251 => x"c3",
          7252 => x"80",
          7253 => x"2e",
          7254 => x"9a",
          7255 => x"7a",
          7256 => x"dd",
          7257 => x"84",
          7258 => x"9d",
          7259 => x"0a",
          7260 => x"51",
          7261 => x"ff",
          7262 => x"7d",
          7263 => x"38",
          7264 => x"52",
          7265 => x"9d",
          7266 => x"55",
          7267 => x"62",
          7268 => x"74",
          7269 => x"75",
          7270 => x"7e",
          7271 => x"b2",
          7272 => x"ec",
          7273 => x"38",
          7274 => x"82",
          7275 => x"52",
          7276 => x"9d",
          7277 => x"16",
          7278 => x"56",
          7279 => x"38",
          7280 => x"77",
          7281 => x"8d",
          7282 => x"7d",
          7283 => x"38",
          7284 => x"57",
          7285 => x"83",
          7286 => x"76",
          7287 => x"7a",
          7288 => x"ff",
          7289 => x"82",
          7290 => x"81",
          7291 => x"16",
          7292 => x"56",
          7293 => x"38",
          7294 => x"83",
          7295 => x"86",
          7296 => x"ff",
          7297 => x"38",
          7298 => x"82",
          7299 => x"81",
          7300 => x"06",
          7301 => x"fe",
          7302 => x"53",
          7303 => x"51",
          7304 => x"3f",
          7305 => x"52",
          7306 => x"9b",
          7307 => x"be",
          7308 => x"75",
          7309 => x"81",
          7310 => x"0b",
          7311 => x"77",
          7312 => x"75",
          7313 => x"60",
          7314 => x"80",
          7315 => x"75",
          7316 => x"b6",
          7317 => x"85",
          7318 => x"85",
          7319 => x"2a",
          7320 => x"75",
          7321 => x"82",
          7322 => x"87",
          7323 => x"52",
          7324 => x"51",
          7325 => x"3f",
          7326 => x"ca",
          7327 => x"9b",
          7328 => x"54",
          7329 => x"52",
          7330 => x"97",
          7331 => x"56",
          7332 => x"08",
          7333 => x"53",
          7334 => x"51",
          7335 => x"3f",
          7336 => x"85",
          7337 => x"38",
          7338 => x"56",
          7339 => x"56",
          7340 => x"85",
          7341 => x"75",
          7342 => x"0c",
          7343 => x"04",
          7344 => x"7d",
          7345 => x"80",
          7346 => x"05",
          7347 => x"76",
          7348 => x"38",
          7349 => x"11",
          7350 => x"53",
          7351 => x"79",
          7352 => x"3f",
          7353 => x"09",
          7354 => x"38",
          7355 => x"55",
          7356 => x"db",
          7357 => x"70",
          7358 => x"34",
          7359 => x"74",
          7360 => x"81",
          7361 => x"80",
          7362 => x"55",
          7363 => x"76",
          7364 => x"85",
          7365 => x"3d",
          7366 => x"3d",
          7367 => x"84",
          7368 => x"33",
          7369 => x"8a",
          7370 => x"06",
          7371 => x"52",
          7372 => x"3f",
          7373 => x"56",
          7374 => x"80",
          7375 => x"17",
          7376 => x"8c",
          7377 => x"77",
          7378 => x"16",
          7379 => x"25",
          7380 => x"3d",
          7381 => x"75",
          7382 => x"52",
          7383 => x"cb",
          7384 => x"76",
          7385 => x"81",
          7386 => x"07",
          7387 => x"09",
          7388 => x"51",
          7389 => x"84",
          7390 => x"19",
          7391 => x"8b",
          7392 => x"f9",
          7393 => x"84",
          7394 => x"56",
          7395 => x"a7",
          7396 => x"fc",
          7397 => x"53",
          7398 => x"75",
          7399 => x"80",
          7400 => x"ec",
          7401 => x"84",
          7402 => x"2e",
          7403 => x"87",
          7404 => x"08",
          7405 => x"ff",
          7406 => x"85",
          7407 => x"3d",
          7408 => x"3d",
          7409 => x"80",
          7410 => x"52",
          7411 => x"99",
          7412 => x"74",
          7413 => x"0d",
          7414 => x"0d",
          7415 => x"05",
          7416 => x"86",
          7417 => x"54",
          7418 => x"73",
          7419 => x"fe",
          7420 => x"51",
          7421 => x"98",
          7422 => x"00",
          7423 => x"ff",
          7424 => x"ff",
          7425 => x"ff",
          7426 => x"00",
          7427 => x"8e",
          7428 => x"12",
          7429 => x"19",
          7430 => x"20",
          7431 => x"27",
          7432 => x"2e",
          7433 => x"35",
          7434 => x"3c",
          7435 => x"43",
          7436 => x"4a",
          7437 => x"51",
          7438 => x"58",
          7439 => x"5e",
          7440 => x"64",
          7441 => x"6a",
          7442 => x"70",
          7443 => x"76",
          7444 => x"7c",
          7445 => x"82",
          7446 => x"88",
          7447 => x"ce",
          7448 => x"d4",
          7449 => x"da",
          7450 => x"e0",
          7451 => x"e6",
          7452 => x"e6",
          7453 => x"d0",
          7454 => x"bd",
          7455 => x"eb",
          7456 => x"b8",
          7457 => x"c3",
          7458 => x"67",
          7459 => x"c2",
          7460 => x"a4",
          7461 => x"3b",
          7462 => x"c0",
          7463 => x"6d",
          7464 => x"c3",
          7465 => x"bd",
          7466 => x"e0",
          7467 => x"67",
          7468 => x"c3",
          7469 => x"c3",
          7470 => x"c0",
          7471 => x"3b",
          7472 => x"c2",
          7473 => x"eb",
          7474 => x"69",
          7475 => x"00",
          7476 => x"63",
          7477 => x"00",
          7478 => x"69",
          7479 => x"00",
          7480 => x"61",
          7481 => x"00",
          7482 => x"65",
          7483 => x"00",
          7484 => x"65",
          7485 => x"00",
          7486 => x"70",
          7487 => x"00",
          7488 => x"66",
          7489 => x"00",
          7490 => x"6d",
          7491 => x"00",
          7492 => x"00",
          7493 => x"00",
          7494 => x"00",
          7495 => x"00",
          7496 => x"00",
          7497 => x"00",
          7498 => x"00",
          7499 => x"6c",
          7500 => x"00",
          7501 => x"00",
          7502 => x"74",
          7503 => x"00",
          7504 => x"65",
          7505 => x"00",
          7506 => x"6f",
          7507 => x"00",
          7508 => x"74",
          7509 => x"00",
          7510 => x"73",
          7511 => x"00",
          7512 => x"73",
          7513 => x"00",
          7514 => x"6f",
          7515 => x"00",
          7516 => x"00",
          7517 => x"6b",
          7518 => x"72",
          7519 => x"00",
          7520 => x"65",
          7521 => x"6c",
          7522 => x"72",
          7523 => x"0a",
          7524 => x"00",
          7525 => x"6b",
          7526 => x"74",
          7527 => x"61",
          7528 => x"0a",
          7529 => x"00",
          7530 => x"66",
          7531 => x"20",
          7532 => x"6e",
          7533 => x"00",
          7534 => x"70",
          7535 => x"20",
          7536 => x"6e",
          7537 => x"00",
          7538 => x"61",
          7539 => x"20",
          7540 => x"65",
          7541 => x"65",
          7542 => x"00",
          7543 => x"65",
          7544 => x"64",
          7545 => x"65",
          7546 => x"00",
          7547 => x"65",
          7548 => x"72",
          7549 => x"79",
          7550 => x"69",
          7551 => x"2e",
          7552 => x"00",
          7553 => x"65",
          7554 => x"6e",
          7555 => x"20",
          7556 => x"61",
          7557 => x"2e",
          7558 => x"00",
          7559 => x"69",
          7560 => x"72",
          7561 => x"20",
          7562 => x"74",
          7563 => x"65",
          7564 => x"00",
          7565 => x"76",
          7566 => x"75",
          7567 => x"72",
          7568 => x"20",
          7569 => x"61",
          7570 => x"2e",
          7571 => x"00",
          7572 => x"6b",
          7573 => x"74",
          7574 => x"61",
          7575 => x"64",
          7576 => x"00",
          7577 => x"63",
          7578 => x"61",
          7579 => x"6c",
          7580 => x"69",
          7581 => x"79",
          7582 => x"6d",
          7583 => x"75",
          7584 => x"6f",
          7585 => x"69",
          7586 => x"0a",
          7587 => x"00",
          7588 => x"6d",
          7589 => x"61",
          7590 => x"74",
          7591 => x"0a",
          7592 => x"00",
          7593 => x"65",
          7594 => x"2c",
          7595 => x"65",
          7596 => x"69",
          7597 => x"63",
          7598 => x"65",
          7599 => x"64",
          7600 => x"00",
          7601 => x"65",
          7602 => x"20",
          7603 => x"6b",
          7604 => x"0a",
          7605 => x"00",
          7606 => x"75",
          7607 => x"63",
          7608 => x"74",
          7609 => x"6d",
          7610 => x"2e",
          7611 => x"00",
          7612 => x"20",
          7613 => x"79",
          7614 => x"65",
          7615 => x"69",
          7616 => x"2e",
          7617 => x"00",
          7618 => x"61",
          7619 => x"65",
          7620 => x"69",
          7621 => x"72",
          7622 => x"74",
          7623 => x"00",
          7624 => x"63",
          7625 => x"2e",
          7626 => x"00",
          7627 => x"6e",
          7628 => x"20",
          7629 => x"6f",
          7630 => x"00",
          7631 => x"75",
          7632 => x"74",
          7633 => x"25",
          7634 => x"74",
          7635 => x"75",
          7636 => x"74",
          7637 => x"73",
          7638 => x"0a",
          7639 => x"00",
          7640 => x"64",
          7641 => x"00",
          7642 => x"58",
          7643 => x"00",
          7644 => x"00",
          7645 => x"58",
          7646 => x"00",
          7647 => x"20",
          7648 => x"20",
          7649 => x"00",
          7650 => x"58",
          7651 => x"00",
          7652 => x"00",
          7653 => x"00",
          7654 => x"00",
          7655 => x"00",
          7656 => x"20",
          7657 => x"28",
          7658 => x"00",
          7659 => x"30",
          7660 => x"30",
          7661 => x"00",
          7662 => x"30",
          7663 => x"00",
          7664 => x"55",
          7665 => x"65",
          7666 => x"30",
          7667 => x"20",
          7668 => x"25",
          7669 => x"2a",
          7670 => x"00",
          7671 => x"20",
          7672 => x"65",
          7673 => x"70",
          7674 => x"61",
          7675 => x"65",
          7676 => x"00",
          7677 => x"65",
          7678 => x"6e",
          7679 => x"72",
          7680 => x"0a",
          7681 => x"00",
          7682 => x"20",
          7683 => x"65",
          7684 => x"70",
          7685 => x"00",
          7686 => x"54",
          7687 => x"44",
          7688 => x"74",
          7689 => x"75",
          7690 => x"00",
          7691 => x"54",
          7692 => x"52",
          7693 => x"74",
          7694 => x"75",
          7695 => x"00",
          7696 => x"54",
          7697 => x"58",
          7698 => x"74",
          7699 => x"75",
          7700 => x"00",
          7701 => x"54",
          7702 => x"58",
          7703 => x"74",
          7704 => x"75",
          7705 => x"00",
          7706 => x"54",
          7707 => x"58",
          7708 => x"74",
          7709 => x"75",
          7710 => x"00",
          7711 => x"54",
          7712 => x"58",
          7713 => x"74",
          7714 => x"75",
          7715 => x"00",
          7716 => x"74",
          7717 => x"20",
          7718 => x"74",
          7719 => x"72",
          7720 => x"0a",
          7721 => x"00",
          7722 => x"62",
          7723 => x"67",
          7724 => x"6d",
          7725 => x"2e",
          7726 => x"00",
          7727 => x"6f",
          7728 => x"63",
          7729 => x"74",
          7730 => x"00",
          7731 => x"2e",
          7732 => x"00",
          7733 => x"00",
          7734 => x"6c",
          7735 => x"74",
          7736 => x"6e",
          7737 => x"61",
          7738 => x"65",
          7739 => x"20",
          7740 => x"64",
          7741 => x"20",
          7742 => x"61",
          7743 => x"69",
          7744 => x"20",
          7745 => x"75",
          7746 => x"79",
          7747 => x"00",
          7748 => x"00",
          7749 => x"61",
          7750 => x"67",
          7751 => x"2e",
          7752 => x"00",
          7753 => x"79",
          7754 => x"2e",
          7755 => x"00",
          7756 => x"70",
          7757 => x"6e",
          7758 => x"2e",
          7759 => x"00",
          7760 => x"6c",
          7761 => x"30",
          7762 => x"2d",
          7763 => x"38",
          7764 => x"25",
          7765 => x"29",
          7766 => x"00",
          7767 => x"70",
          7768 => x"6d",
          7769 => x"0a",
          7770 => x"00",
          7771 => x"6d",
          7772 => x"74",
          7773 => x"00",
          7774 => x"58",
          7775 => x"32",
          7776 => x"00",
          7777 => x"0a",
          7778 => x"00",
          7779 => x"58",
          7780 => x"34",
          7781 => x"00",
          7782 => x"58",
          7783 => x"38",
          7784 => x"00",
          7785 => x"63",
          7786 => x"6e",
          7787 => x"6f",
          7788 => x"40",
          7789 => x"38",
          7790 => x"2e",
          7791 => x"00",
          7792 => x"6c",
          7793 => x"20",
          7794 => x"65",
          7795 => x"25",
          7796 => x"20",
          7797 => x"0a",
          7798 => x"00",
          7799 => x"6c",
          7800 => x"74",
          7801 => x"65",
          7802 => x"6f",
          7803 => x"28",
          7804 => x"2e",
          7805 => x"00",
          7806 => x"74",
          7807 => x"69",
          7808 => x"61",
          7809 => x"69",
          7810 => x"69",
          7811 => x"2e",
          7812 => x"00",
          7813 => x"64",
          7814 => x"62",
          7815 => x"69",
          7816 => x"2e",
          7817 => x"00",
          7818 => x"00",
          7819 => x"00",
          7820 => x"5c",
          7821 => x"25",
          7822 => x"73",
          7823 => x"00",
          7824 => x"5c",
          7825 => x"25",
          7826 => x"00",
          7827 => x"5c",
          7828 => x"00",
          7829 => x"20",
          7830 => x"6d",
          7831 => x"2e",
          7832 => x"00",
          7833 => x"6e",
          7834 => x"2e",
          7835 => x"00",
          7836 => x"62",
          7837 => x"67",
          7838 => x"74",
          7839 => x"75",
          7840 => x"2e",
          7841 => x"00",
          7842 => x"25",
          7843 => x"64",
          7844 => x"3a",
          7845 => x"25",
          7846 => x"64",
          7847 => x"00",
          7848 => x"20",
          7849 => x"66",
          7850 => x"72",
          7851 => x"6f",
          7852 => x"00",
          7853 => x"72",
          7854 => x"53",
          7855 => x"63",
          7856 => x"69",
          7857 => x"00",
          7858 => x"65",
          7859 => x"65",
          7860 => x"6d",
          7861 => x"6d",
          7862 => x"65",
          7863 => x"00",
          7864 => x"20",
          7865 => x"53",
          7866 => x"4d",
          7867 => x"25",
          7868 => x"3a",
          7869 => x"58",
          7870 => x"00",
          7871 => x"20",
          7872 => x"41",
          7873 => x"20",
          7874 => x"25",
          7875 => x"3a",
          7876 => x"58",
          7877 => x"00",
          7878 => x"20",
          7879 => x"4e",
          7880 => x"41",
          7881 => x"25",
          7882 => x"3a",
          7883 => x"58",
          7884 => x"00",
          7885 => x"20",
          7886 => x"4d",
          7887 => x"20",
          7888 => x"25",
          7889 => x"3a",
          7890 => x"58",
          7891 => x"00",
          7892 => x"20",
          7893 => x"20",
          7894 => x"20",
          7895 => x"25",
          7896 => x"3a",
          7897 => x"58",
          7898 => x"00",
          7899 => x"20",
          7900 => x"43",
          7901 => x"20",
          7902 => x"44",
          7903 => x"63",
          7904 => x"3d",
          7905 => x"64",
          7906 => x"00",
          7907 => x"20",
          7908 => x"45",
          7909 => x"20",
          7910 => x"54",
          7911 => x"72",
          7912 => x"3d",
          7913 => x"64",
          7914 => x"00",
          7915 => x"20",
          7916 => x"52",
          7917 => x"52",
          7918 => x"43",
          7919 => x"6e",
          7920 => x"3d",
          7921 => x"64",
          7922 => x"00",
          7923 => x"20",
          7924 => x"48",
          7925 => x"45",
          7926 => x"53",
          7927 => x"00",
          7928 => x"20",
          7929 => x"49",
          7930 => x"00",
          7931 => x"20",
          7932 => x"54",
          7933 => x"00",
          7934 => x"20",
          7935 => x"0a",
          7936 => x"00",
          7937 => x"20",
          7938 => x"0a",
          7939 => x"00",
          7940 => x"72",
          7941 => x"65",
          7942 => x"00",
          7943 => x"20",
          7944 => x"20",
          7945 => x"65",
          7946 => x"65",
          7947 => x"72",
          7948 => x"64",
          7949 => x"73",
          7950 => x"25",
          7951 => x"0a",
          7952 => x"00",
          7953 => x"20",
          7954 => x"20",
          7955 => x"6f",
          7956 => x"53",
          7957 => x"74",
          7958 => x"64",
          7959 => x"73",
          7960 => x"25",
          7961 => x"0a",
          7962 => x"00",
          7963 => x"20",
          7964 => x"63",
          7965 => x"74",
          7966 => x"20",
          7967 => x"72",
          7968 => x"20",
          7969 => x"20",
          7970 => x"25",
          7971 => x"0a",
          7972 => x"00",
          7973 => x"63",
          7974 => x"00",
          7975 => x"20",
          7976 => x"20",
          7977 => x"20",
          7978 => x"20",
          7979 => x"20",
          7980 => x"20",
          7981 => x"20",
          7982 => x"25",
          7983 => x"0a",
          7984 => x"00",
          7985 => x"20",
          7986 => x"74",
          7987 => x"43",
          7988 => x"6b",
          7989 => x"65",
          7990 => x"20",
          7991 => x"20",
          7992 => x"25",
          7993 => x"30",
          7994 => x"48",
          7995 => x"00",
          7996 => x"20",
          7997 => x"41",
          7998 => x"6c",
          7999 => x"20",
          8000 => x"71",
          8001 => x"20",
          8002 => x"20",
          8003 => x"25",
          8004 => x"30",
          8005 => x"48",
          8006 => x"00",
          8007 => x"20",
          8008 => x"68",
          8009 => x"65",
          8010 => x"52",
          8011 => x"43",
          8012 => x"6b",
          8013 => x"65",
          8014 => x"25",
          8015 => x"30",
          8016 => x"48",
          8017 => x"00",
          8018 => x"6c",
          8019 => x"00",
          8020 => x"69",
          8021 => x"00",
          8022 => x"78",
          8023 => x"00",
          8024 => x"00",
          8025 => x"6d",
          8026 => x"00",
          8027 => x"6e",
          8028 => x"00",
          8029 => x"d0",
          8030 => x"00",
          8031 => x"02",
          8032 => x"cc",
          8033 => x"00",
          8034 => x"03",
          8035 => x"c8",
          8036 => x"00",
          8037 => x"04",
          8038 => x"c4",
          8039 => x"00",
          8040 => x"05",
          8041 => x"c0",
          8042 => x"00",
          8043 => x"06",
          8044 => x"bc",
          8045 => x"00",
          8046 => x"07",
          8047 => x"b8",
          8048 => x"00",
          8049 => x"01",
          8050 => x"b4",
          8051 => x"00",
          8052 => x"08",
          8053 => x"b0",
          8054 => x"00",
          8055 => x"0b",
          8056 => x"ac",
          8057 => x"00",
          8058 => x"09",
          8059 => x"a8",
          8060 => x"00",
          8061 => x"0a",
          8062 => x"a4",
          8063 => x"00",
          8064 => x"0d",
          8065 => x"a0",
          8066 => x"00",
          8067 => x"0c",
          8068 => x"9c",
          8069 => x"00",
          8070 => x"0e",
          8071 => x"98",
          8072 => x"00",
          8073 => x"0f",
          8074 => x"94",
          8075 => x"00",
          8076 => x"0f",
          8077 => x"90",
          8078 => x"00",
          8079 => x"10",
          8080 => x"8c",
          8081 => x"00",
          8082 => x"11",
          8083 => x"88",
          8084 => x"00",
          8085 => x"12",
          8086 => x"84",
          8087 => x"00",
          8088 => x"13",
          8089 => x"80",
          8090 => x"00",
          8091 => x"14",
          8092 => x"7c",
          8093 => x"00",
          8094 => x"15",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"7e",
          8100 => x"7e",
          8101 => x"7e",
          8102 => x"00",
          8103 => x"7e",
          8104 => x"7e",
          8105 => x"7e",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"74",
          8118 => x"00",
          8119 => x"74",
          8120 => x"00",
          8121 => x"00",
          8122 => x"64",
          8123 => x"73",
          8124 => x"00",
          8125 => x"6c",
          8126 => x"74",
          8127 => x"65",
          8128 => x"20",
          8129 => x"20",
          8130 => x"74",
          8131 => x"20",
          8132 => x"65",
          8133 => x"20",
          8134 => x"2e",
          8135 => x"00",
          8136 => x"6e",
          8137 => x"6f",
          8138 => x"2f",
          8139 => x"61",
          8140 => x"68",
          8141 => x"6f",
          8142 => x"66",
          8143 => x"2c",
          8144 => x"73",
          8145 => x"69",
          8146 => x"0a",
          8147 => x"00",
          8148 => x"00",
          8149 => x"2c",
          8150 => x"3d",
          8151 => x"5d",
          8152 => x"00",
          8153 => x"00",
          8154 => x"33",
          8155 => x"00",
          8156 => x"4d",
          8157 => x"53",
          8158 => x"00",
          8159 => x"4e",
          8160 => x"20",
          8161 => x"46",
          8162 => x"32",
          8163 => x"00",
          8164 => x"4e",
          8165 => x"20",
          8166 => x"46",
          8167 => x"20",
          8168 => x"00",
          8169 => x"50",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"41",
          8174 => x"80",
          8175 => x"49",
          8176 => x"8f",
          8177 => x"4f",
          8178 => x"55",
          8179 => x"9b",
          8180 => x"9f",
          8181 => x"55",
          8182 => x"a7",
          8183 => x"ab",
          8184 => x"af",
          8185 => x"b3",
          8186 => x"b7",
          8187 => x"bb",
          8188 => x"bf",
          8189 => x"c3",
          8190 => x"c7",
          8191 => x"cb",
          8192 => x"cf",
          8193 => x"d3",
          8194 => x"d7",
          8195 => x"db",
          8196 => x"df",
          8197 => x"e3",
          8198 => x"e7",
          8199 => x"eb",
          8200 => x"ef",
          8201 => x"f3",
          8202 => x"f7",
          8203 => x"fb",
          8204 => x"ff",
          8205 => x"3b",
          8206 => x"2f",
          8207 => x"3a",
          8208 => x"7c",
          8209 => x"00",
          8210 => x"04",
          8211 => x"40",
          8212 => x"00",
          8213 => x"00",
          8214 => x"02",
          8215 => x"08",
          8216 => x"20",
          8217 => x"00",
          8218 => x"00",
          8219 => x"c8",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"d0",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"d8",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"e0",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"e8",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"f0",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"f8",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"08",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"10",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"14",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"18",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"1c",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"20",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"24",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"28",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"2c",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"34",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"38",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"40",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"48",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"50",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"58",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"60",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"68",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"70",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"ff",
          8326 => x"00",
          8327 => x"ff",
          8328 => x"00",
          8329 => x"ff",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"ff",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"01",
          8343 => x"01",
          8344 => x"01",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"d4",
          8371 => x"00",
          8372 => x"dc",
          8373 => x"00",
          8374 => x"e4",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"83",
             1 => x"0b",
             2 => x"9b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"92",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"81",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a5",
           270 => x"0b",
           271 => x"0b",
           272 => x"c5",
           273 => x"0b",
           274 => x"0b",
           275 => x"e5",
           276 => x"0b",
           277 => x"0b",
           278 => x"85",
           279 => x"0b",
           280 => x"0b",
           281 => x"a5",
           282 => x"0b",
           283 => x"0b",
           284 => x"c5",
           285 => x"0b",
           286 => x"0b",
           287 => x"e5",
           288 => x"0b",
           289 => x"0b",
           290 => x"84",
           291 => x"0b",
           292 => x"0b",
           293 => x"a2",
           294 => x"0b",
           295 => x"0b",
           296 => x"c2",
           297 => x"0b",
           298 => x"0b",
           299 => x"e2",
           300 => x"0b",
           301 => x"0b",
           302 => x"82",
           303 => x"0b",
           304 => x"0b",
           305 => x"a2",
           306 => x"0b",
           307 => x"0b",
           308 => x"c2",
           309 => x"0b",
           310 => x"0b",
           311 => x"e2",
           312 => x"0b",
           313 => x"0b",
           314 => x"82",
           315 => x"0b",
           316 => x"0b",
           317 => x"a2",
           318 => x"0b",
           319 => x"0b",
           320 => x"c2",
           321 => x"0b",
           322 => x"0b",
           323 => x"e2",
           324 => x"0b",
           325 => x"0b",
           326 => x"82",
           327 => x"0b",
           328 => x"0b",
           329 => x"a2",
           330 => x"0b",
           331 => x"0b",
           332 => x"c2",
           333 => x"0b",
           334 => x"0b",
           335 => x"e2",
           336 => x"0b",
           337 => x"0b",
           338 => x"82",
           339 => x"0b",
           340 => x"0b",
           341 => x"a0",
           342 => x"0b",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"85",
           386 => x"c1",
           387 => x"85",
           388 => x"a0",
           389 => x"85",
           390 => x"ce",
           391 => x"85",
           392 => x"a0",
           393 => x"85",
           394 => x"ce",
           395 => x"85",
           396 => x"a0",
           397 => x"85",
           398 => x"ce",
           399 => x"85",
           400 => x"a0",
           401 => x"85",
           402 => x"d5",
           403 => x"85",
           404 => x"a0",
           405 => x"85",
           406 => x"d6",
           407 => x"85",
           408 => x"a0",
           409 => x"85",
           410 => x"cf",
           411 => x"85",
           412 => x"a0",
           413 => x"85",
           414 => x"d6",
           415 => x"85",
           416 => x"a0",
           417 => x"85",
           418 => x"d8",
           419 => x"85",
           420 => x"a0",
           421 => x"85",
           422 => x"d4",
           423 => x"85",
           424 => x"a0",
           425 => x"85",
           426 => x"cf",
           427 => x"85",
           428 => x"a0",
           429 => x"85",
           430 => x"d4",
           431 => x"85",
           432 => x"a0",
           433 => x"85",
           434 => x"d5",
           435 => x"85",
           436 => x"a0",
           437 => x"85",
           438 => x"c3",
           439 => x"85",
           440 => x"a0",
           441 => x"85",
           442 => x"c3",
           443 => x"85",
           444 => x"a0",
           445 => x"85",
           446 => x"c4",
           447 => x"f8",
           448 => x"90",
           449 => x"f8",
           450 => x"2d",
           451 => x"08",
           452 => x"04",
           453 => x"0c",
           454 => x"82",
           455 => x"82",
           456 => x"82",
           457 => x"81",
           458 => x"82",
           459 => x"82",
           460 => x"82",
           461 => x"81",
           462 => x"82",
           463 => x"82",
           464 => x"82",
           465 => x"81",
           466 => x"82",
           467 => x"82",
           468 => x"82",
           469 => x"81",
           470 => x"82",
           471 => x"82",
           472 => x"82",
           473 => x"81",
           474 => x"82",
           475 => x"82",
           476 => x"82",
           477 => x"81",
           478 => x"82",
           479 => x"82",
           480 => x"82",
           481 => x"81",
           482 => x"82",
           483 => x"82",
           484 => x"82",
           485 => x"81",
           486 => x"82",
           487 => x"82",
           488 => x"82",
           489 => x"81",
           490 => x"82",
           491 => x"82",
           492 => x"82",
           493 => x"81",
           494 => x"82",
           495 => x"82",
           496 => x"82",
           497 => x"81",
           498 => x"82",
           499 => x"82",
           500 => x"82",
           501 => x"81",
           502 => x"82",
           503 => x"82",
           504 => x"82",
           505 => x"81",
           506 => x"82",
           507 => x"82",
           508 => x"82",
           509 => x"81",
           510 => x"82",
           511 => x"82",
           512 => x"82",
           513 => x"81",
           514 => x"82",
           515 => x"82",
           516 => x"82",
           517 => x"81",
           518 => x"82",
           519 => x"82",
           520 => x"82",
           521 => x"81",
           522 => x"82",
           523 => x"82",
           524 => x"82",
           525 => x"81",
           526 => x"82",
           527 => x"82",
           528 => x"82",
           529 => x"81",
           530 => x"82",
           531 => x"82",
           532 => x"82",
           533 => x"81",
           534 => x"82",
           535 => x"82",
           536 => x"82",
           537 => x"81",
           538 => x"82",
           539 => x"82",
           540 => x"82",
           541 => x"81",
           542 => x"82",
           543 => x"82",
           544 => x"82",
           545 => x"81",
           546 => x"82",
           547 => x"82",
           548 => x"82",
           549 => x"81",
           550 => x"82",
           551 => x"82",
           552 => x"82",
           553 => x"81",
           554 => x"82",
           555 => x"82",
           556 => x"82",
           557 => x"81",
           558 => x"82",
           559 => x"82",
           560 => x"82",
           561 => x"81",
           562 => x"82",
           563 => x"82",
           564 => x"82",
           565 => x"80",
           566 => x"82",
           567 => x"82",
           568 => x"82",
           569 => x"80",
           570 => x"82",
           571 => x"82",
           572 => x"82",
           573 => x"80",
           574 => x"82",
           575 => x"82",
           576 => x"82",
           577 => x"bb",
           578 => x"85",
           579 => x"a0",
           580 => x"85",
           581 => x"93",
           582 => x"f8",
           583 => x"90",
           584 => x"f8",
           585 => x"80",
           586 => x"f8",
           587 => x"90",
           588 => x"f8",
           589 => x"2d",
           590 => x"08",
           591 => x"04",
           592 => x"00",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"10",
           598 => x"10",
           599 => x"10",
           600 => x"53",
           601 => x"00",
           602 => x"06",
           603 => x"09",
           604 => x"05",
           605 => x"2b",
           606 => x"06",
           607 => x"04",
           608 => x"72",
           609 => x"05",
           610 => x"05",
           611 => x"72",
           612 => x"53",
           613 => x"51",
           614 => x"04",
           615 => x"70",
           616 => x"27",
           617 => x"71",
           618 => x"53",
           619 => x"0b",
           620 => x"8c",
           621 => x"9d",
           622 => x"85",
           623 => x"82",
           624 => x"fe",
           625 => x"85",
           626 => x"05",
           627 => x"f8",
           628 => x"0c",
           629 => x"08",
           630 => x"52",
           631 => x"85",
           632 => x"05",
           633 => x"82",
           634 => x"fc",
           635 => x"81",
           636 => x"51",
           637 => x"83",
           638 => x"82",
           639 => x"fc",
           640 => x"05",
           641 => x"08",
           642 => x"82",
           643 => x"fc",
           644 => x"85",
           645 => x"05",
           646 => x"82",
           647 => x"51",
           648 => x"82",
           649 => x"04",
           650 => x"08",
           651 => x"f8",
           652 => x"0d",
           653 => x"08",
           654 => x"82",
           655 => x"fc",
           656 => x"85",
           657 => x"05",
           658 => x"33",
           659 => x"08",
           660 => x"81",
           661 => x"f8",
           662 => x"0c",
           663 => x"08",
           664 => x"53",
           665 => x"34",
           666 => x"08",
           667 => x"81",
           668 => x"f8",
           669 => x"0c",
           670 => x"06",
           671 => x"2e",
           672 => x"be",
           673 => x"f8",
           674 => x"08",
           675 => x"ec",
           676 => x"3d",
           677 => x"f8",
           678 => x"85",
           679 => x"82",
           680 => x"fd",
           681 => x"85",
           682 => x"05",
           683 => x"f8",
           684 => x"0c",
           685 => x"08",
           686 => x"82",
           687 => x"f8",
           688 => x"85",
           689 => x"05",
           690 => x"80",
           691 => x"85",
           692 => x"05",
           693 => x"82",
           694 => x"90",
           695 => x"85",
           696 => x"05",
           697 => x"82",
           698 => x"90",
           699 => x"85",
           700 => x"05",
           701 => x"ba",
           702 => x"f8",
           703 => x"08",
           704 => x"82",
           705 => x"f8",
           706 => x"05",
           707 => x"08",
           708 => x"82",
           709 => x"fc",
           710 => x"52",
           711 => x"82",
           712 => x"fc",
           713 => x"05",
           714 => x"08",
           715 => x"ff",
           716 => x"85",
           717 => x"05",
           718 => x"85",
           719 => x"85",
           720 => x"85",
           721 => x"82",
           722 => x"02",
           723 => x"0c",
           724 => x"82",
           725 => x"90",
           726 => x"2e",
           727 => x"82",
           728 => x"8c",
           729 => x"71",
           730 => x"f8",
           731 => x"08",
           732 => x"85",
           733 => x"05",
           734 => x"f8",
           735 => x"08",
           736 => x"81",
           737 => x"54",
           738 => x"71",
           739 => x"80",
           740 => x"85",
           741 => x"05",
           742 => x"33",
           743 => x"08",
           744 => x"81",
           745 => x"f8",
           746 => x"0c",
           747 => x"06",
           748 => x"8d",
           749 => x"82",
           750 => x"fc",
           751 => x"9b",
           752 => x"f8",
           753 => x"08",
           754 => x"85",
           755 => x"05",
           756 => x"f8",
           757 => x"08",
           758 => x"38",
           759 => x"82",
           760 => x"90",
           761 => x"2e",
           762 => x"82",
           763 => x"88",
           764 => x"33",
           765 => x"8d",
           766 => x"82",
           767 => x"fc",
           768 => x"d7",
           769 => x"f8",
           770 => x"08",
           771 => x"85",
           772 => x"05",
           773 => x"f8",
           774 => x"08",
           775 => x"52",
           776 => x"81",
           777 => x"f8",
           778 => x"0c",
           779 => x"85",
           780 => x"05",
           781 => x"82",
           782 => x"8c",
           783 => x"33",
           784 => x"70",
           785 => x"08",
           786 => x"53",
           787 => x"53",
           788 => x"0b",
           789 => x"08",
           790 => x"82",
           791 => x"fc",
           792 => x"85",
           793 => x"3d",
           794 => x"f8",
           795 => x"85",
           796 => x"82",
           797 => x"fe",
           798 => x"85",
           799 => x"05",
           800 => x"f8",
           801 => x"0c",
           802 => x"08",
           803 => x"80",
           804 => x"38",
           805 => x"08",
           806 => x"81",
           807 => x"f8",
           808 => x"0c",
           809 => x"08",
           810 => x"ff",
           811 => x"f8",
           812 => x"0c",
           813 => x"08",
           814 => x"80",
           815 => x"82",
           816 => x"8c",
           817 => x"70",
           818 => x"08",
           819 => x"52",
           820 => x"34",
           821 => x"08",
           822 => x"81",
           823 => x"f8",
           824 => x"0c",
           825 => x"82",
           826 => x"88",
           827 => x"82",
           828 => x"51",
           829 => x"82",
           830 => x"04",
           831 => x"08",
           832 => x"f8",
           833 => x"0d",
           834 => x"85",
           835 => x"05",
           836 => x"f8",
           837 => x"08",
           838 => x"38",
           839 => x"08",
           840 => x"30",
           841 => x"08",
           842 => x"80",
           843 => x"f8",
           844 => x"0c",
           845 => x"08",
           846 => x"8a",
           847 => x"82",
           848 => x"f4",
           849 => x"85",
           850 => x"05",
           851 => x"f8",
           852 => x"0c",
           853 => x"08",
           854 => x"80",
           855 => x"82",
           856 => x"8c",
           857 => x"82",
           858 => x"8c",
           859 => x"0b",
           860 => x"08",
           861 => x"82",
           862 => x"fc",
           863 => x"38",
           864 => x"85",
           865 => x"05",
           866 => x"f8",
           867 => x"08",
           868 => x"08",
           869 => x"80",
           870 => x"f8",
           871 => x"08",
           872 => x"f8",
           873 => x"08",
           874 => x"3f",
           875 => x"08",
           876 => x"f8",
           877 => x"0c",
           878 => x"f8",
           879 => x"08",
           880 => x"38",
           881 => x"08",
           882 => x"30",
           883 => x"08",
           884 => x"82",
           885 => x"f8",
           886 => x"82",
           887 => x"54",
           888 => x"82",
           889 => x"04",
           890 => x"08",
           891 => x"f8",
           892 => x"0d",
           893 => x"85",
           894 => x"05",
           895 => x"f8",
           896 => x"08",
           897 => x"38",
           898 => x"08",
           899 => x"30",
           900 => x"08",
           901 => x"81",
           902 => x"f8",
           903 => x"0c",
           904 => x"08",
           905 => x"80",
           906 => x"82",
           907 => x"8c",
           908 => x"82",
           909 => x"8c",
           910 => x"53",
           911 => x"08",
           912 => x"52",
           913 => x"08",
           914 => x"51",
           915 => x"82",
           916 => x"70",
           917 => x"08",
           918 => x"54",
           919 => x"08",
           920 => x"80",
           921 => x"82",
           922 => x"f8",
           923 => x"82",
           924 => x"f8",
           925 => x"85",
           926 => x"05",
           927 => x"85",
           928 => x"87",
           929 => x"85",
           930 => x"82",
           931 => x"02",
           932 => x"0c",
           933 => x"80",
           934 => x"f8",
           935 => x"0c",
           936 => x"08",
           937 => x"81",
           938 => x"70",
           939 => x"85",
           940 => x"05",
           941 => x"85",
           942 => x"05",
           943 => x"85",
           944 => x"05",
           945 => x"f8",
           946 => x"08",
           947 => x"85",
           948 => x"05",
           949 => x"f8",
           950 => x"08",
           951 => x"f8",
           952 => x"0c",
           953 => x"51",
           954 => x"08",
           955 => x"80",
           956 => x"ff",
           957 => x"85",
           958 => x"05",
           959 => x"85",
           960 => x"83",
           961 => x"85",
           962 => x"82",
           963 => x"02",
           964 => x"0c",
           965 => x"80",
           966 => x"f8",
           967 => x"08",
           968 => x"f8",
           969 => x"08",
           970 => x"3f",
           971 => x"08",
           972 => x"ec",
           973 => x"3d",
           974 => x"f8",
           975 => x"85",
           976 => x"82",
           977 => x"fd",
           978 => x"53",
           979 => x"08",
           980 => x"52",
           981 => x"08",
           982 => x"51",
           983 => x"85",
           984 => x"82",
           985 => x"54",
           986 => x"82",
           987 => x"04",
           988 => x"08",
           989 => x"f8",
           990 => x"0d",
           991 => x"85",
           992 => x"05",
           993 => x"82",
           994 => x"f8",
           995 => x"85",
           996 => x"05",
           997 => x"f8",
           998 => x"08",
           999 => x"82",
          1000 => x"fc",
          1001 => x"2e",
          1002 => x"0b",
          1003 => x"08",
          1004 => x"24",
          1005 => x"85",
          1006 => x"05",
          1007 => x"85",
          1008 => x"05",
          1009 => x"f8",
          1010 => x"08",
          1011 => x"f8",
          1012 => x"0c",
          1013 => x"82",
          1014 => x"fc",
          1015 => x"2e",
          1016 => x"82",
          1017 => x"8c",
          1018 => x"85",
          1019 => x"05",
          1020 => x"38",
          1021 => x"08",
          1022 => x"82",
          1023 => x"8c",
          1024 => x"82",
          1025 => x"88",
          1026 => x"85",
          1027 => x"05",
          1028 => x"f8",
          1029 => x"08",
          1030 => x"f8",
          1031 => x"0c",
          1032 => x"08",
          1033 => x"81",
          1034 => x"f8",
          1035 => x"0c",
          1036 => x"08",
          1037 => x"81",
          1038 => x"f8",
          1039 => x"0c",
          1040 => x"82",
          1041 => x"90",
          1042 => x"2e",
          1043 => x"85",
          1044 => x"05",
          1045 => x"85",
          1046 => x"05",
          1047 => x"39",
          1048 => x"08",
          1049 => x"70",
          1050 => x"08",
          1051 => x"51",
          1052 => x"08",
          1053 => x"82",
          1054 => x"85",
          1055 => x"85",
          1056 => x"f9",
          1057 => x"70",
          1058 => x"56",
          1059 => x"2e",
          1060 => x"95",
          1061 => x"51",
          1062 => x"82",
          1063 => x"15",
          1064 => x"16",
          1065 => x"cd",
          1066 => x"54",
          1067 => x"09",
          1068 => x"38",
          1069 => x"f1",
          1070 => x"76",
          1071 => x"80",
          1072 => x"08",
          1073 => x"f2",
          1074 => x"ec",
          1075 => x"52",
          1076 => x"f4",
          1077 => x"85",
          1078 => x"38",
          1079 => x"54",
          1080 => x"ff",
          1081 => x"17",
          1082 => x"06",
          1083 => x"77",
          1084 => x"ff",
          1085 => x"85",
          1086 => x"3d",
          1087 => x"3d",
          1088 => x"71",
          1089 => x"8d",
          1090 => x"2b",
          1091 => x"8c",
          1092 => x"81",
          1093 => x"81",
          1094 => x"eb",
          1095 => x"f9",
          1096 => x"94",
          1097 => x"39",
          1098 => x"51",
          1099 => x"81",
          1100 => x"80",
          1101 => x"eb",
          1102 => x"dd",
          1103 => x"dc",
          1104 => x"39",
          1105 => x"51",
          1106 => x"81",
          1107 => x"80",
          1108 => x"ec",
          1109 => x"c1",
          1110 => x"b4",
          1111 => x"81",
          1112 => x"b5",
          1113 => x"e4",
          1114 => x"81",
          1115 => x"a9",
          1116 => x"a4",
          1117 => x"81",
          1118 => x"9d",
          1119 => x"d8",
          1120 => x"81",
          1121 => x"91",
          1122 => x"88",
          1123 => x"81",
          1124 => x"85",
          1125 => x"ac",
          1126 => x"3f",
          1127 => x"04",
          1128 => x"77",
          1129 => x"74",
          1130 => x"92",
          1131 => x"52",
          1132 => x"d7",
          1133 => x"82",
          1134 => x"51",
          1135 => x"e8",
          1136 => x"fa",
          1137 => x"85",
          1138 => x"75",
          1139 => x"3f",
          1140 => x"08",
          1141 => x"75",
          1142 => x"bc",
          1143 => x"3f",
          1144 => x"04",
          1145 => x"66",
          1146 => x"80",
          1147 => x"5b",
          1148 => x"78",
          1149 => x"70",
          1150 => x"25",
          1151 => x"59",
          1152 => x"87",
          1153 => x"38",
          1154 => x"76",
          1155 => x"ff",
          1156 => x"93",
          1157 => x"86",
          1158 => x"76",
          1159 => x"70",
          1160 => x"86",
          1161 => x"85",
          1162 => x"82",
          1163 => x"b9",
          1164 => x"ec",
          1165 => x"98",
          1166 => x"85",
          1167 => x"96",
          1168 => x"54",
          1169 => x"77",
          1170 => x"81",
          1171 => x"82",
          1172 => x"57",
          1173 => x"08",
          1174 => x"55",
          1175 => x"89",
          1176 => x"75",
          1177 => x"d7",
          1178 => x"d8",
          1179 => x"92",
          1180 => x"09",
          1181 => x"78",
          1182 => x"7b",
          1183 => x"70",
          1184 => x"06",
          1185 => x"56",
          1186 => x"90",
          1187 => x"e0",
          1188 => x"98",
          1189 => x"78",
          1190 => x"3f",
          1191 => x"82",
          1192 => x"96",
          1193 => x"f9",
          1194 => x"02",
          1195 => x"05",
          1196 => x"ff",
          1197 => x"7a",
          1198 => x"fe",
          1199 => x"85",
          1200 => x"38",
          1201 => x"88",
          1202 => x"2e",
          1203 => x"39",
          1204 => x"54",
          1205 => x"53",
          1206 => x"51",
          1207 => x"85",
          1208 => x"83",
          1209 => x"76",
          1210 => x"0c",
          1211 => x"04",
          1212 => x"7f",
          1213 => x"8c",
          1214 => x"05",
          1215 => x"15",
          1216 => x"5c",
          1217 => x"5e",
          1218 => x"ee",
          1219 => x"cc",
          1220 => x"f0",
          1221 => x"3f",
          1222 => x"79",
          1223 => x"38",
          1224 => x"89",
          1225 => x"2e",
          1226 => x"c1",
          1227 => x"53",
          1228 => x"8d",
          1229 => x"52",
          1230 => x"51",
          1231 => x"88",
          1232 => x"80",
          1233 => x"3f",
          1234 => x"bf",
          1235 => x"53",
          1236 => x"8d",
          1237 => x"52",
          1238 => x"51",
          1239 => x"88",
          1240 => x"fc",
          1241 => x"3f",
          1242 => x"9f",
          1243 => x"53",
          1244 => x"8d",
          1245 => x"52",
          1246 => x"51",
          1247 => x"88",
          1248 => x"90",
          1249 => x"3f",
          1250 => x"a0",
          1251 => x"3f",
          1252 => x"81",
          1253 => x"a7",
          1254 => x"55",
          1255 => x"bb",
          1256 => x"70",
          1257 => x"80",
          1258 => x"27",
          1259 => x"56",
          1260 => x"74",
          1261 => x"81",
          1262 => x"06",
          1263 => x"06",
          1264 => x"80",
          1265 => x"73",
          1266 => x"85",
          1267 => x"83",
          1268 => x"a6",
          1269 => x"15",
          1270 => x"81",
          1271 => x"a7",
          1272 => x"18",
          1273 => x"58",
          1274 => x"82",
          1275 => x"98",
          1276 => x"2c",
          1277 => x"a0",
          1278 => x"06",
          1279 => x"e5",
          1280 => x"ec",
          1281 => x"70",
          1282 => x"a0",
          1283 => x"81",
          1284 => x"32",
          1285 => x"05",
          1286 => x"73",
          1287 => x"51",
          1288 => x"57",
          1289 => x"73",
          1290 => x"76",
          1291 => x"81",
          1292 => x"80",
          1293 => x"7c",
          1294 => x"78",
          1295 => x"38",
          1296 => x"82",
          1297 => x"8f",
          1298 => x"fc",
          1299 => x"9b",
          1300 => x"ef",
          1301 => x"ef",
          1302 => x"ab",
          1303 => x"84",
          1304 => x"a4",
          1305 => x"ef",
          1306 => x"ef",
          1307 => x"84",
          1308 => x"81",
          1309 => x"ab",
          1310 => x"80",
          1311 => x"a0",
          1312 => x"3d",
          1313 => x"3d",
          1314 => x"96",
          1315 => x"a4",
          1316 => x"51",
          1317 => x"81",
          1318 => x"98",
          1319 => x"51",
          1320 => x"72",
          1321 => x"81",
          1322 => x"71",
          1323 => x"38",
          1324 => x"cd",
          1325 => x"f4",
          1326 => x"3f",
          1327 => x"c1",
          1328 => x"2a",
          1329 => x"51",
          1330 => x"2e",
          1331 => x"51",
          1332 => x"81",
          1333 => x"98",
          1334 => x"51",
          1335 => x"72",
          1336 => x"81",
          1337 => x"71",
          1338 => x"38",
          1339 => x"91",
          1340 => x"98",
          1341 => x"3f",
          1342 => x"85",
          1343 => x"2a",
          1344 => x"51",
          1345 => x"2e",
          1346 => x"51",
          1347 => x"81",
          1348 => x"97",
          1349 => x"51",
          1350 => x"72",
          1351 => x"81",
          1352 => x"71",
          1353 => x"38",
          1354 => x"d5",
          1355 => x"c0",
          1356 => x"3f",
          1357 => x"c9",
          1358 => x"2a",
          1359 => x"51",
          1360 => x"2e",
          1361 => x"51",
          1362 => x"81",
          1363 => x"97",
          1364 => x"51",
          1365 => x"72",
          1366 => x"81",
          1367 => x"71",
          1368 => x"38",
          1369 => x"99",
          1370 => x"e8",
          1371 => x"3f",
          1372 => x"8d",
          1373 => x"2a",
          1374 => x"51",
          1375 => x"2e",
          1376 => x"51",
          1377 => x"81",
          1378 => x"96",
          1379 => x"51",
          1380 => x"a2",
          1381 => x"3d",
          1382 => x"3d",
          1383 => x"84",
          1384 => x"33",
          1385 => x"56",
          1386 => x"51",
          1387 => x"0b",
          1388 => x"e8",
          1389 => x"ab",
          1390 => x"81",
          1391 => x"82",
          1392 => x"80",
          1393 => x"82",
          1394 => x"09",
          1395 => x"82",
          1396 => x"07",
          1397 => x"71",
          1398 => x"54",
          1399 => x"82",
          1400 => x"0b",
          1401 => x"e8",
          1402 => x"81",
          1403 => x"06",
          1404 => x"9c",
          1405 => x"52",
          1406 => x"b9",
          1407 => x"85",
          1408 => x"2e",
          1409 => x"85",
          1410 => x"a2",
          1411 => x"39",
          1412 => x"51",
          1413 => x"3f",
          1414 => x"0b",
          1415 => x"34",
          1416 => x"80",
          1417 => x"73",
          1418 => x"81",
          1419 => x"81",
          1420 => x"74",
          1421 => x"b5",
          1422 => x"0b",
          1423 => x"0c",
          1424 => x"04",
          1425 => x"80",
          1426 => x"9c",
          1427 => x"5d",
          1428 => x"51",
          1429 => x"3f",
          1430 => x"08",
          1431 => x"59",
          1432 => x"09",
          1433 => x"38",
          1434 => x"52",
          1435 => x"52",
          1436 => x"3f",
          1437 => x"52",
          1438 => x"51",
          1439 => x"3f",
          1440 => x"08",
          1441 => x"38",
          1442 => x"51",
          1443 => x"81",
          1444 => x"81",
          1445 => x"a1",
          1446 => x"3d",
          1447 => x"80",
          1448 => x"51",
          1449 => x"b4",
          1450 => x"05",
          1451 => x"3f",
          1452 => x"08",
          1453 => x"90",
          1454 => x"78",
          1455 => x"87",
          1456 => x"80",
          1457 => x"38",
          1458 => x"81",
          1459 => x"bd",
          1460 => x"78",
          1461 => x"bb",
          1462 => x"2e",
          1463 => x"8a",
          1464 => x"80",
          1465 => x"94",
          1466 => x"c0",
          1467 => x"38",
          1468 => x"82",
          1469 => x"a4",
          1470 => x"f9",
          1471 => x"38",
          1472 => x"24",
          1473 => x"80",
          1474 => x"fa",
          1475 => x"f8",
          1476 => x"38",
          1477 => x"78",
          1478 => x"89",
          1479 => x"81",
          1480 => x"38",
          1481 => x"2e",
          1482 => x"89",
          1483 => x"81",
          1484 => x"e2",
          1485 => x"39",
          1486 => x"80",
          1487 => x"84",
          1488 => x"90",
          1489 => x"ec",
          1490 => x"fe",
          1491 => x"3d",
          1492 => x"53",
          1493 => x"51",
          1494 => x"82",
          1495 => x"80",
          1496 => x"38",
          1497 => x"f8",
          1498 => x"84",
          1499 => x"e4",
          1500 => x"ec",
          1501 => x"82",
          1502 => x"42",
          1503 => x"51",
          1504 => x"63",
          1505 => x"79",
          1506 => x"e9",
          1507 => x"78",
          1508 => x"05",
          1509 => x"7a",
          1510 => x"81",
          1511 => x"3d",
          1512 => x"53",
          1513 => x"51",
          1514 => x"82",
          1515 => x"80",
          1516 => x"38",
          1517 => x"fc",
          1518 => x"84",
          1519 => x"94",
          1520 => x"ec",
          1521 => x"fd",
          1522 => x"3d",
          1523 => x"53",
          1524 => x"51",
          1525 => x"82",
          1526 => x"80",
          1527 => x"38",
          1528 => x"51",
          1529 => x"63",
          1530 => x"27",
          1531 => x"61",
          1532 => x"81",
          1533 => x"79",
          1534 => x"05",
          1535 => x"b4",
          1536 => x"11",
          1537 => x"05",
          1538 => x"3f",
          1539 => x"08",
          1540 => x"ff",
          1541 => x"fe",
          1542 => x"ff",
          1543 => x"a6",
          1544 => x"85",
          1545 => x"2e",
          1546 => x"b4",
          1547 => x"11",
          1548 => x"05",
          1549 => x"3f",
          1550 => x"08",
          1551 => x"d3",
          1552 => x"b0",
          1553 => x"3f",
          1554 => x"63",
          1555 => x"61",
          1556 => x"33",
          1557 => x"78",
          1558 => x"38",
          1559 => x"54",
          1560 => x"79",
          1561 => x"c0",
          1562 => x"3f",
          1563 => x"81",
          1564 => x"d6",
          1565 => x"d8",
          1566 => x"39",
          1567 => x"80",
          1568 => x"84",
          1569 => x"cc",
          1570 => x"ec",
          1571 => x"38",
          1572 => x"33",
          1573 => x"2e",
          1574 => x"84",
          1575 => x"80",
          1576 => x"84",
          1577 => x"78",
          1578 => x"38",
          1579 => x"08",
          1580 => x"82",
          1581 => x"59",
          1582 => x"88",
          1583 => x"a0",
          1584 => x"39",
          1585 => x"33",
          1586 => x"2e",
          1587 => x"84",
          1588 => x"9a",
          1589 => x"d6",
          1590 => x"80",
          1591 => x"82",
          1592 => x"44",
          1593 => x"84",
          1594 => x"80",
          1595 => x"3d",
          1596 => x"53",
          1597 => x"51",
          1598 => x"82",
          1599 => x"80",
          1600 => x"84",
          1601 => x"78",
          1602 => x"38",
          1603 => x"08",
          1604 => x"39",
          1605 => x"33",
          1606 => x"2e",
          1607 => x"84",
          1608 => x"bb",
          1609 => x"da",
          1610 => x"80",
          1611 => x"82",
          1612 => x"43",
          1613 => x"84",
          1614 => x"78",
          1615 => x"38",
          1616 => x"08",
          1617 => x"82",
          1618 => x"59",
          1619 => x"88",
          1620 => x"b4",
          1621 => x"39",
          1622 => x"08",
          1623 => x"b4",
          1624 => x"11",
          1625 => x"05",
          1626 => x"3f",
          1627 => x"08",
          1628 => x"38",
          1629 => x"5c",
          1630 => x"83",
          1631 => x"7a",
          1632 => x"09",
          1633 => x"72",
          1634 => x"70",
          1635 => x"51",
          1636 => x"80",
          1637 => x"7a",
          1638 => x"38",
          1639 => x"f2",
          1640 => x"c8",
          1641 => x"63",
          1642 => x"62",
          1643 => x"f2",
          1644 => x"f2",
          1645 => x"b4",
          1646 => x"39",
          1647 => x"80",
          1648 => x"84",
          1649 => x"8c",
          1650 => x"ec",
          1651 => x"f9",
          1652 => x"3d",
          1653 => x"53",
          1654 => x"51",
          1655 => x"82",
          1656 => x"80",
          1657 => x"63",
          1658 => x"cb",
          1659 => x"34",
          1660 => x"44",
          1661 => x"fc",
          1662 => x"84",
          1663 => x"d4",
          1664 => x"ec",
          1665 => x"f9",
          1666 => x"70",
          1667 => x"81",
          1668 => x"a0",
          1669 => x"f8",
          1670 => x"a1",
          1671 => x"45",
          1672 => x"78",
          1673 => x"eb",
          1674 => x"27",
          1675 => x"3d",
          1676 => x"53",
          1677 => x"51",
          1678 => x"82",
          1679 => x"80",
          1680 => x"63",
          1681 => x"cb",
          1682 => x"34",
          1683 => x"44",
          1684 => x"81",
          1685 => x"9a",
          1686 => x"ae",
          1687 => x"fe",
          1688 => x"ff",
          1689 => x"a3",
          1690 => x"85",
          1691 => x"2e",
          1692 => x"b4",
          1693 => x"11",
          1694 => x"05",
          1695 => x"3f",
          1696 => x"08",
          1697 => x"38",
          1698 => x"be",
          1699 => x"70",
          1700 => x"23",
          1701 => x"3d",
          1702 => x"53",
          1703 => x"51",
          1704 => x"82",
          1705 => x"e0",
          1706 => x"39",
          1707 => x"54",
          1708 => x"8c",
          1709 => x"3f",
          1710 => x"79",
          1711 => x"3f",
          1712 => x"33",
          1713 => x"2e",
          1714 => x"78",
          1715 => x"38",
          1716 => x"41",
          1717 => x"3d",
          1718 => x"53",
          1719 => x"51",
          1720 => x"82",
          1721 => x"80",
          1722 => x"60",
          1723 => x"05",
          1724 => x"82",
          1725 => x"78",
          1726 => x"39",
          1727 => x"51",
          1728 => x"ff",
          1729 => x"3d",
          1730 => x"53",
          1731 => x"51",
          1732 => x"82",
          1733 => x"80",
          1734 => x"38",
          1735 => x"f0",
          1736 => x"84",
          1737 => x"a8",
          1738 => x"ec",
          1739 => x"a0",
          1740 => x"71",
          1741 => x"84",
          1742 => x"3d",
          1743 => x"53",
          1744 => x"51",
          1745 => x"82",
          1746 => x"e5",
          1747 => x"39",
          1748 => x"54",
          1749 => x"98",
          1750 => x"3f",
          1751 => x"79",
          1752 => x"3f",
          1753 => x"33",
          1754 => x"2e",
          1755 => x"9f",
          1756 => x"38",
          1757 => x"f0",
          1758 => x"84",
          1759 => x"d0",
          1760 => x"ec",
          1761 => x"8d",
          1762 => x"71",
          1763 => x"84",
          1764 => x"bc",
          1765 => x"84",
          1766 => x"3f",
          1767 => x"b4",
          1768 => x"11",
          1769 => x"05",
          1770 => x"3f",
          1771 => x"08",
          1772 => x"df",
          1773 => x"81",
          1774 => x"9d",
          1775 => x"59",
          1776 => x"3d",
          1777 => x"53",
          1778 => x"51",
          1779 => x"82",
          1780 => x"80",
          1781 => x"38",
          1782 => x"f3",
          1783 => x"fc",
          1784 => x"78",
          1785 => x"ec",
          1786 => x"f5",
          1787 => x"85",
          1788 => x"81",
          1789 => x"9c",
          1790 => x"97",
          1791 => x"f8",
          1792 => x"3f",
          1793 => x"f5",
          1794 => x"f4",
          1795 => x"dc",
          1796 => x"ff",
          1797 => x"ef",
          1798 => x"39",
          1799 => x"33",
          1800 => x"2e",
          1801 => x"7d",
          1802 => x"78",
          1803 => x"d0",
          1804 => x"ff",
          1805 => x"83",
          1806 => x"85",
          1807 => x"81",
          1808 => x"2e",
          1809 => x"82",
          1810 => x"7a",
          1811 => x"38",
          1812 => x"7a",
          1813 => x"38",
          1814 => x"81",
          1815 => x"7b",
          1816 => x"ac",
          1817 => x"81",
          1818 => x"b4",
          1819 => x"05",
          1820 => x"3f",
          1821 => x"f4",
          1822 => x"3d",
          1823 => x"51",
          1824 => x"a9",
          1825 => x"81",
          1826 => x"80",
          1827 => x"c0",
          1828 => x"ff",
          1829 => x"9b",
          1830 => x"39",
          1831 => x"53",
          1832 => x"52",
          1833 => x"b0",
          1834 => x"c6",
          1835 => x"90",
          1836 => x"fc",
          1837 => x"64",
          1838 => x"82",
          1839 => x"82",
          1840 => x"b4",
          1841 => x"05",
          1842 => x"3f",
          1843 => x"08",
          1844 => x"08",
          1845 => x"81",
          1846 => x"07",
          1847 => x"5b",
          1848 => x"5a",
          1849 => x"83",
          1850 => x"78",
          1851 => x"78",
          1852 => x"38",
          1853 => x"81",
          1854 => x"59",
          1855 => x"38",
          1856 => x"7d",
          1857 => x"59",
          1858 => x"7e",
          1859 => x"81",
          1860 => x"38",
          1861 => x"51",
          1862 => x"f2",
          1863 => x"3d",
          1864 => x"82",
          1865 => x"87",
          1866 => x"70",
          1867 => x"87",
          1868 => x"72",
          1869 => x"3f",
          1870 => x"08",
          1871 => x"08",
          1872 => x"84",
          1873 => x"51",
          1874 => x"72",
          1875 => x"08",
          1876 => x"87",
          1877 => x"70",
          1878 => x"87",
          1879 => x"72",
          1880 => x"3f",
          1881 => x"08",
          1882 => x"08",
          1883 => x"84",
          1884 => x"51",
          1885 => x"72",
          1886 => x"08",
          1887 => x"8c",
          1888 => x"87",
          1889 => x"0c",
          1890 => x"0b",
          1891 => x"94",
          1892 => x"9a",
          1893 => x"f4",
          1894 => x"95",
          1895 => x"f8",
          1896 => x"3f",
          1897 => x"81",
          1898 => x"93",
          1899 => x"f4",
          1900 => x"b8",
          1901 => x"51",
          1902 => x"81",
          1903 => x"3f",
          1904 => x"80",
          1905 => x"0d",
          1906 => x"53",
          1907 => x"52",
          1908 => x"82",
          1909 => x"81",
          1910 => x"07",
          1911 => x"52",
          1912 => x"e8",
          1913 => x"85",
          1914 => x"3d",
          1915 => x"3d",
          1916 => x"08",
          1917 => x"73",
          1918 => x"74",
          1919 => x"38",
          1920 => x"70",
          1921 => x"81",
          1922 => x"81",
          1923 => x"39",
          1924 => x"70",
          1925 => x"81",
          1926 => x"81",
          1927 => x"54",
          1928 => x"81",
          1929 => x"06",
          1930 => x"39",
          1931 => x"80",
          1932 => x"54",
          1933 => x"83",
          1934 => x"70",
          1935 => x"38",
          1936 => x"98",
          1937 => x"52",
          1938 => x"52",
          1939 => x"2e",
          1940 => x"54",
          1941 => x"84",
          1942 => x"38",
          1943 => x"52",
          1944 => x"2e",
          1945 => x"83",
          1946 => x"70",
          1947 => x"09",
          1948 => x"80",
          1949 => x"51",
          1950 => x"80",
          1951 => x"80",
          1952 => x"05",
          1953 => x"75",
          1954 => x"70",
          1955 => x"0c",
          1956 => x"04",
          1957 => x"76",
          1958 => x"80",
          1959 => x"86",
          1960 => x"52",
          1961 => x"a8",
          1962 => x"ec",
          1963 => x"80",
          1964 => x"74",
          1965 => x"85",
          1966 => x"3d",
          1967 => x"3d",
          1968 => x"11",
          1969 => x"52",
          1970 => x"70",
          1971 => x"98",
          1972 => x"33",
          1973 => x"82",
          1974 => x"26",
          1975 => x"84",
          1976 => x"83",
          1977 => x"26",
          1978 => x"85",
          1979 => x"84",
          1980 => x"26",
          1981 => x"86",
          1982 => x"85",
          1983 => x"26",
          1984 => x"88",
          1985 => x"86",
          1986 => x"e7",
          1987 => x"38",
          1988 => x"54",
          1989 => x"87",
          1990 => x"cc",
          1991 => x"87",
          1992 => x"0c",
          1993 => x"c0",
          1994 => x"82",
          1995 => x"c0",
          1996 => x"83",
          1997 => x"c0",
          1998 => x"84",
          1999 => x"c0",
          2000 => x"85",
          2001 => x"c0",
          2002 => x"86",
          2003 => x"c0",
          2004 => x"74",
          2005 => x"a4",
          2006 => x"c0",
          2007 => x"80",
          2008 => x"98",
          2009 => x"52",
          2010 => x"ec",
          2011 => x"0d",
          2012 => x"0d",
          2013 => x"c0",
          2014 => x"81",
          2015 => x"c0",
          2016 => x"5e",
          2017 => x"87",
          2018 => x"08",
          2019 => x"1c",
          2020 => x"98",
          2021 => x"79",
          2022 => x"87",
          2023 => x"08",
          2024 => x"1c",
          2025 => x"98",
          2026 => x"79",
          2027 => x"87",
          2028 => x"08",
          2029 => x"1c",
          2030 => x"98",
          2031 => x"7b",
          2032 => x"87",
          2033 => x"08",
          2034 => x"1c",
          2035 => x"0c",
          2036 => x"ff",
          2037 => x"83",
          2038 => x"58",
          2039 => x"57",
          2040 => x"56",
          2041 => x"55",
          2042 => x"54",
          2043 => x"53",
          2044 => x"ff",
          2045 => x"f5",
          2046 => x"e0",
          2047 => x"0d",
          2048 => x"0d",
          2049 => x"33",
          2050 => x"05",
          2051 => x"51",
          2052 => x"82",
          2053 => x"83",
          2054 => x"fb",
          2055 => x"82",
          2056 => x"70",
          2057 => x"57",
          2058 => x"c0",
          2059 => x"74",
          2060 => x"38",
          2061 => x"94",
          2062 => x"70",
          2063 => x"81",
          2064 => x"52",
          2065 => x"8c",
          2066 => x"2a",
          2067 => x"51",
          2068 => x"38",
          2069 => x"70",
          2070 => x"51",
          2071 => x"8d",
          2072 => x"2a",
          2073 => x"51",
          2074 => x"be",
          2075 => x"ff",
          2076 => x"c0",
          2077 => x"70",
          2078 => x"38",
          2079 => x"90",
          2080 => x"0c",
          2081 => x"ec",
          2082 => x"0d",
          2083 => x"0d",
          2084 => x"33",
          2085 => x"33",
          2086 => x"06",
          2087 => x"87",
          2088 => x"51",
          2089 => x"86",
          2090 => x"94",
          2091 => x"08",
          2092 => x"70",
          2093 => x"54",
          2094 => x"2e",
          2095 => x"91",
          2096 => x"06",
          2097 => x"d7",
          2098 => x"32",
          2099 => x"51",
          2100 => x"2e",
          2101 => x"93",
          2102 => x"06",
          2103 => x"ff",
          2104 => x"81",
          2105 => x"87",
          2106 => x"52",
          2107 => x"86",
          2108 => x"94",
          2109 => x"72",
          2110 => x"0d",
          2111 => x"0d",
          2112 => x"74",
          2113 => x"ff",
          2114 => x"57",
          2115 => x"80",
          2116 => x"81",
          2117 => x"15",
          2118 => x"33",
          2119 => x"06",
          2120 => x"58",
          2121 => x"84",
          2122 => x"2e",
          2123 => x"c0",
          2124 => x"70",
          2125 => x"2a",
          2126 => x"53",
          2127 => x"80",
          2128 => x"71",
          2129 => x"81",
          2130 => x"70",
          2131 => x"81",
          2132 => x"06",
          2133 => x"80",
          2134 => x"71",
          2135 => x"81",
          2136 => x"70",
          2137 => x"74",
          2138 => x"51",
          2139 => x"80",
          2140 => x"2e",
          2141 => x"c0",
          2142 => x"77",
          2143 => x"17",
          2144 => x"81",
          2145 => x"53",
          2146 => x"86",
          2147 => x"85",
          2148 => x"3d",
          2149 => x"3d",
          2150 => x"8c",
          2151 => x"ff",
          2152 => x"87",
          2153 => x"51",
          2154 => x"86",
          2155 => x"94",
          2156 => x"08",
          2157 => x"70",
          2158 => x"51",
          2159 => x"2e",
          2160 => x"81",
          2161 => x"87",
          2162 => x"52",
          2163 => x"86",
          2164 => x"94",
          2165 => x"08",
          2166 => x"06",
          2167 => x"0c",
          2168 => x"0d",
          2169 => x"0d",
          2170 => x"33",
          2171 => x"06",
          2172 => x"c0",
          2173 => x"70",
          2174 => x"38",
          2175 => x"94",
          2176 => x"70",
          2177 => x"81",
          2178 => x"51",
          2179 => x"80",
          2180 => x"72",
          2181 => x"51",
          2182 => x"80",
          2183 => x"2e",
          2184 => x"c0",
          2185 => x"71",
          2186 => x"2b",
          2187 => x"51",
          2188 => x"82",
          2189 => x"84",
          2190 => x"ff",
          2191 => x"c0",
          2192 => x"70",
          2193 => x"06",
          2194 => x"80",
          2195 => x"38",
          2196 => x"a4",
          2197 => x"90",
          2198 => x"9e",
          2199 => x"84",
          2200 => x"c0",
          2201 => x"82",
          2202 => x"87",
          2203 => x"08",
          2204 => x"0c",
          2205 => x"9c",
          2206 => x"a0",
          2207 => x"9e",
          2208 => x"84",
          2209 => x"c0",
          2210 => x"82",
          2211 => x"87",
          2212 => x"08",
          2213 => x"0c",
          2214 => x"b4",
          2215 => x"b0",
          2216 => x"9e",
          2217 => x"84",
          2218 => x"c0",
          2219 => x"82",
          2220 => x"87",
          2221 => x"08",
          2222 => x"0c",
          2223 => x"c4",
          2224 => x"c0",
          2225 => x"9e",
          2226 => x"70",
          2227 => x"23",
          2228 => x"84",
          2229 => x"c8",
          2230 => x"9e",
          2231 => x"84",
          2232 => x"c0",
          2233 => x"82",
          2234 => x"81",
          2235 => x"d4",
          2236 => x"87",
          2237 => x"08",
          2238 => x"0a",
          2239 => x"52",
          2240 => x"83",
          2241 => x"71",
          2242 => x"34",
          2243 => x"c0",
          2244 => x"70",
          2245 => x"06",
          2246 => x"70",
          2247 => x"38",
          2248 => x"82",
          2249 => x"80",
          2250 => x"9e",
          2251 => x"90",
          2252 => x"51",
          2253 => x"80",
          2254 => x"81",
          2255 => x"84",
          2256 => x"0b",
          2257 => x"90",
          2258 => x"80",
          2259 => x"52",
          2260 => x"2e",
          2261 => x"52",
          2262 => x"d8",
          2263 => x"87",
          2264 => x"08",
          2265 => x"80",
          2266 => x"52",
          2267 => x"83",
          2268 => x"71",
          2269 => x"34",
          2270 => x"c0",
          2271 => x"70",
          2272 => x"06",
          2273 => x"70",
          2274 => x"38",
          2275 => x"82",
          2276 => x"80",
          2277 => x"9e",
          2278 => x"84",
          2279 => x"51",
          2280 => x"80",
          2281 => x"81",
          2282 => x"84",
          2283 => x"0b",
          2284 => x"90",
          2285 => x"80",
          2286 => x"52",
          2287 => x"2e",
          2288 => x"52",
          2289 => x"dc",
          2290 => x"87",
          2291 => x"08",
          2292 => x"80",
          2293 => x"52",
          2294 => x"83",
          2295 => x"71",
          2296 => x"34",
          2297 => x"c0",
          2298 => x"70",
          2299 => x"06",
          2300 => x"70",
          2301 => x"38",
          2302 => x"82",
          2303 => x"80",
          2304 => x"9e",
          2305 => x"a0",
          2306 => x"52",
          2307 => x"2e",
          2308 => x"52",
          2309 => x"df",
          2310 => x"9e",
          2311 => x"98",
          2312 => x"8a",
          2313 => x"51",
          2314 => x"e0",
          2315 => x"87",
          2316 => x"08",
          2317 => x"06",
          2318 => x"70",
          2319 => x"38",
          2320 => x"82",
          2321 => x"87",
          2322 => x"08",
          2323 => x"06",
          2324 => x"51",
          2325 => x"82",
          2326 => x"80",
          2327 => x"9e",
          2328 => x"88",
          2329 => x"52",
          2330 => x"83",
          2331 => x"71",
          2332 => x"34",
          2333 => x"90",
          2334 => x"06",
          2335 => x"82",
          2336 => x"83",
          2337 => x"fc",
          2338 => x"f5",
          2339 => x"dc",
          2340 => x"d4",
          2341 => x"80",
          2342 => x"81",
          2343 => x"85",
          2344 => x"f5",
          2345 => x"c4",
          2346 => x"d6",
          2347 => x"80",
          2348 => x"82",
          2349 => x"82",
          2350 => x"11",
          2351 => x"f5",
          2352 => x"98",
          2353 => x"db",
          2354 => x"80",
          2355 => x"82",
          2356 => x"82",
          2357 => x"11",
          2358 => x"f5",
          2359 => x"fc",
          2360 => x"d8",
          2361 => x"80",
          2362 => x"82",
          2363 => x"82",
          2364 => x"11",
          2365 => x"f6",
          2366 => x"e0",
          2367 => x"d9",
          2368 => x"80",
          2369 => x"82",
          2370 => x"82",
          2371 => x"11",
          2372 => x"f6",
          2373 => x"c4",
          2374 => x"da",
          2375 => x"80",
          2376 => x"82",
          2377 => x"82",
          2378 => x"11",
          2379 => x"f6",
          2380 => x"a8",
          2381 => x"df",
          2382 => x"80",
          2383 => x"82",
          2384 => x"52",
          2385 => x"51",
          2386 => x"82",
          2387 => x"54",
          2388 => x"8d",
          2389 => x"e4",
          2390 => x"f7",
          2391 => x"fc",
          2392 => x"e1",
          2393 => x"80",
          2394 => x"82",
          2395 => x"52",
          2396 => x"51",
          2397 => x"82",
          2398 => x"54",
          2399 => x"88",
          2400 => x"cc",
          2401 => x"3f",
          2402 => x"33",
          2403 => x"2e",
          2404 => x"f7",
          2405 => x"d4",
          2406 => x"dc",
          2407 => x"80",
          2408 => x"81",
          2409 => x"83",
          2410 => x"84",
          2411 => x"73",
          2412 => x"38",
          2413 => x"51",
          2414 => x"82",
          2415 => x"54",
          2416 => x"88",
          2417 => x"84",
          2418 => x"3f",
          2419 => x"51",
          2420 => x"82",
          2421 => x"52",
          2422 => x"51",
          2423 => x"82",
          2424 => x"52",
          2425 => x"51",
          2426 => x"82",
          2427 => x"52",
          2428 => x"51",
          2429 => x"81",
          2430 => x"82",
          2431 => x"84",
          2432 => x"81",
          2433 => x"88",
          2434 => x"84",
          2435 => x"bd",
          2436 => x"74",
          2437 => x"3f",
          2438 => x"08",
          2439 => x"c0",
          2440 => x"ec",
          2441 => x"e3",
          2442 => x"85",
          2443 => x"53",
          2444 => x"f9",
          2445 => x"a4",
          2446 => x"db",
          2447 => x"80",
          2448 => x"82",
          2449 => x"55",
          2450 => x"52",
          2451 => x"bb",
          2452 => x"ec",
          2453 => x"84",
          2454 => x"85",
          2455 => x"d0",
          2456 => x"82",
          2457 => x"31",
          2458 => x"81",
          2459 => x"87",
          2460 => x"84",
          2461 => x"73",
          2462 => x"38",
          2463 => x"08",
          2464 => x"c0",
          2465 => x"d1",
          2466 => x"85",
          2467 => x"bd",
          2468 => x"82",
          2469 => x"51",
          2470 => x"74",
          2471 => x"08",
          2472 => x"52",
          2473 => x"51",
          2474 => x"81",
          2475 => x"81",
          2476 => x"3d",
          2477 => x"3d",
          2478 => x"05",
          2479 => x"52",
          2480 => x"a9",
          2481 => x"2b",
          2482 => x"dc",
          2483 => x"81",
          2484 => x"9d",
          2485 => x"d0",
          2486 => x"81",
          2487 => x"91",
          2488 => x"e0",
          2489 => x"81",
          2490 => x"85",
          2491 => x"ec",
          2492 => x"3f",
          2493 => x"04",
          2494 => x"0c",
          2495 => x"87",
          2496 => x"0c",
          2497 => x"e8",
          2498 => x"96",
          2499 => x"fe",
          2500 => x"93",
          2501 => x"72",
          2502 => x"81",
          2503 => x"8d",
          2504 => x"82",
          2505 => x"52",
          2506 => x"90",
          2507 => x"34",
          2508 => x"08",
          2509 => x"9c",
          2510 => x"39",
          2511 => x"08",
          2512 => x"2e",
          2513 => x"51",
          2514 => x"3d",
          2515 => x"3d",
          2516 => x"05",
          2517 => x"f4",
          2518 => x"9c",
          2519 => x"51",
          2520 => x"72",
          2521 => x"0c",
          2522 => x"04",
          2523 => x"75",
          2524 => x"70",
          2525 => x"53",
          2526 => x"2e",
          2527 => x"81",
          2528 => x"81",
          2529 => x"87",
          2530 => x"85",
          2531 => x"fc",
          2532 => x"82",
          2533 => x"78",
          2534 => x"0c",
          2535 => x"33",
          2536 => x"06",
          2537 => x"80",
          2538 => x"72",
          2539 => x"51",
          2540 => x"fe",
          2541 => x"39",
          2542 => x"f4",
          2543 => x"0d",
          2544 => x"0d",
          2545 => x"59",
          2546 => x"05",
          2547 => x"75",
          2548 => x"84",
          2549 => x"2e",
          2550 => x"82",
          2551 => x"70",
          2552 => x"05",
          2553 => x"5b",
          2554 => x"2e",
          2555 => x"85",
          2556 => x"8b",
          2557 => x"2e",
          2558 => x"8a",
          2559 => x"78",
          2560 => x"5a",
          2561 => x"aa",
          2562 => x"06",
          2563 => x"84",
          2564 => x"7b",
          2565 => x"5d",
          2566 => x"59",
          2567 => x"d0",
          2568 => x"89",
          2569 => x"7a",
          2570 => x"11",
          2571 => x"d0",
          2572 => x"81",
          2573 => x"59",
          2574 => x"e3",
          2575 => x"ec",
          2576 => x"81",
          2577 => x"07",
          2578 => x"80",
          2579 => x"09",
          2580 => x"72",
          2581 => x"73",
          2582 => x"58",
          2583 => x"73",
          2584 => x"38",
          2585 => x"79",
          2586 => x"5b",
          2587 => x"75",
          2588 => x"e4",
          2589 => x"80",
          2590 => x"89",
          2591 => x"70",
          2592 => x"55",
          2593 => x"cf",
          2594 => x"38",
          2595 => x"24",
          2596 => x"80",
          2597 => x"8e",
          2598 => x"c3",
          2599 => x"73",
          2600 => x"81",
          2601 => x"99",
          2602 => x"c4",
          2603 => x"38",
          2604 => x"73",
          2605 => x"81",
          2606 => x"80",
          2607 => x"38",
          2608 => x"2e",
          2609 => x"f9",
          2610 => x"d8",
          2611 => x"38",
          2612 => x"77",
          2613 => x"08",
          2614 => x"80",
          2615 => x"55",
          2616 => x"8d",
          2617 => x"70",
          2618 => x"51",
          2619 => x"f5",
          2620 => x"2a",
          2621 => x"74",
          2622 => x"53",
          2623 => x"8f",
          2624 => x"fc",
          2625 => x"81",
          2626 => x"80",
          2627 => x"73",
          2628 => x"3f",
          2629 => x"56",
          2630 => x"27",
          2631 => x"a0",
          2632 => x"3f",
          2633 => x"84",
          2634 => x"33",
          2635 => x"93",
          2636 => x"95",
          2637 => x"91",
          2638 => x"8d",
          2639 => x"89",
          2640 => x"fb",
          2641 => x"80",
          2642 => x"2a",
          2643 => x"51",
          2644 => x"2e",
          2645 => x"84",
          2646 => x"86",
          2647 => x"78",
          2648 => x"08",
          2649 => x"32",
          2650 => x"05",
          2651 => x"80",
          2652 => x"55",
          2653 => x"25",
          2654 => x"80",
          2655 => x"74",
          2656 => x"7a",
          2657 => x"55",
          2658 => x"3d",
          2659 => x"52",
          2660 => x"aa",
          2661 => x"ec",
          2662 => x"06",
          2663 => x"52",
          2664 => x"3f",
          2665 => x"08",
          2666 => x"27",
          2667 => x"14",
          2668 => x"f8",
          2669 => x"87",
          2670 => x"81",
          2671 => x"b0",
          2672 => x"7d",
          2673 => x"5f",
          2674 => x"75",
          2675 => x"70",
          2676 => x"2a",
          2677 => x"76",
          2678 => x"38",
          2679 => x"38",
          2680 => x"70",
          2681 => x"53",
          2682 => x"8e",
          2683 => x"77",
          2684 => x"53",
          2685 => x"81",
          2686 => x"7a",
          2687 => x"55",
          2688 => x"83",
          2689 => x"79",
          2690 => x"81",
          2691 => x"72",
          2692 => x"17",
          2693 => x"27",
          2694 => x"51",
          2695 => x"75",
          2696 => x"72",
          2697 => x"81",
          2698 => x"7a",
          2699 => x"38",
          2700 => x"05",
          2701 => x"ff",
          2702 => x"70",
          2703 => x"57",
          2704 => x"76",
          2705 => x"81",
          2706 => x"72",
          2707 => x"f8",
          2708 => x"f9",
          2709 => x"39",
          2710 => x"04",
          2711 => x"86",
          2712 => x"84",
          2713 => x"55",
          2714 => x"fa",
          2715 => x"3d",
          2716 => x"3d",
          2717 => x"9c",
          2718 => x"3d",
          2719 => x"75",
          2720 => x"3f",
          2721 => x"08",
          2722 => x"34",
          2723 => x"9c",
          2724 => x"3d",
          2725 => x"3d",
          2726 => x"f4",
          2727 => x"9c",
          2728 => x"3d",
          2729 => x"77",
          2730 => x"95",
          2731 => x"9c",
          2732 => x"3d",
          2733 => x"3d",
          2734 => x"82",
          2735 => x"70",
          2736 => x"55",
          2737 => x"80",
          2738 => x"38",
          2739 => x"08",
          2740 => x"82",
          2741 => x"81",
          2742 => x"72",
          2743 => x"ce",
          2744 => x"2e",
          2745 => x"88",
          2746 => x"81",
          2747 => x"25",
          2748 => x"73",
          2749 => x"38",
          2750 => x"86",
          2751 => x"54",
          2752 => x"73",
          2753 => x"ff",
          2754 => x"72",
          2755 => x"38",
          2756 => x"72",
          2757 => x"14",
          2758 => x"f7",
          2759 => x"ac",
          2760 => x"52",
          2761 => x"8a",
          2762 => x"3f",
          2763 => x"82",
          2764 => x"87",
          2765 => x"fe",
          2766 => x"9c",
          2767 => x"82",
          2768 => x"77",
          2769 => x"53",
          2770 => x"72",
          2771 => x"0c",
          2772 => x"04",
          2773 => x"7a",
          2774 => x"80",
          2775 => x"58",
          2776 => x"33",
          2777 => x"a0",
          2778 => x"06",
          2779 => x"13",
          2780 => x"39",
          2781 => x"09",
          2782 => x"38",
          2783 => x"11",
          2784 => x"08",
          2785 => x"54",
          2786 => x"2e",
          2787 => x"80",
          2788 => x"08",
          2789 => x"0c",
          2790 => x"33",
          2791 => x"80",
          2792 => x"38",
          2793 => x"80",
          2794 => x"38",
          2795 => x"57",
          2796 => x"0c",
          2797 => x"33",
          2798 => x"39",
          2799 => x"74",
          2800 => x"38",
          2801 => x"80",
          2802 => x"89",
          2803 => x"38",
          2804 => x"d0",
          2805 => x"55",
          2806 => x"80",
          2807 => x"39",
          2808 => x"e3",
          2809 => x"80",
          2810 => x"27",
          2811 => x"80",
          2812 => x"89",
          2813 => x"70",
          2814 => x"55",
          2815 => x"70",
          2816 => x"55",
          2817 => x"27",
          2818 => x"14",
          2819 => x"06",
          2820 => x"74",
          2821 => x"73",
          2822 => x"38",
          2823 => x"51",
          2824 => x"82",
          2825 => x"14",
          2826 => x"05",
          2827 => x"08",
          2828 => x"54",
          2829 => x"39",
          2830 => x"86",
          2831 => x"81",
          2832 => x"79",
          2833 => x"74",
          2834 => x"0c",
          2835 => x"04",
          2836 => x"7a",
          2837 => x"80",
          2838 => x"58",
          2839 => x"33",
          2840 => x"a0",
          2841 => x"06",
          2842 => x"13",
          2843 => x"39",
          2844 => x"09",
          2845 => x"38",
          2846 => x"11",
          2847 => x"08",
          2848 => x"54",
          2849 => x"2e",
          2850 => x"80",
          2851 => x"08",
          2852 => x"0c",
          2853 => x"33",
          2854 => x"80",
          2855 => x"38",
          2856 => x"80",
          2857 => x"38",
          2858 => x"57",
          2859 => x"0c",
          2860 => x"33",
          2861 => x"39",
          2862 => x"74",
          2863 => x"38",
          2864 => x"80",
          2865 => x"89",
          2866 => x"38",
          2867 => x"d0",
          2868 => x"55",
          2869 => x"80",
          2870 => x"39",
          2871 => x"e3",
          2872 => x"80",
          2873 => x"27",
          2874 => x"80",
          2875 => x"89",
          2876 => x"70",
          2877 => x"55",
          2878 => x"70",
          2879 => x"55",
          2880 => x"27",
          2881 => x"14",
          2882 => x"06",
          2883 => x"74",
          2884 => x"73",
          2885 => x"38",
          2886 => x"51",
          2887 => x"82",
          2888 => x"14",
          2889 => x"05",
          2890 => x"08",
          2891 => x"54",
          2892 => x"39",
          2893 => x"86",
          2894 => x"81",
          2895 => x"79",
          2896 => x"74",
          2897 => x"0c",
          2898 => x"04",
          2899 => x"76",
          2900 => x"98",
          2901 => x"2b",
          2902 => x"72",
          2903 => x"82",
          2904 => x"51",
          2905 => x"80",
          2906 => x"f8",
          2907 => x"52",
          2908 => x"a0",
          2909 => x"fa",
          2910 => x"14",
          2911 => x"97",
          2912 => x"33",
          2913 => x"54",
          2914 => x"09",
          2915 => x"38",
          2916 => x"52",
          2917 => x"ec",
          2918 => x"0d",
          2919 => x"0d",
          2920 => x"05",
          2921 => x"71",
          2922 => x"53",
          2923 => x"9f",
          2924 => x"f2",
          2925 => x"51",
          2926 => x"88",
          2927 => x"3f",
          2928 => x"05",
          2929 => x"34",
          2930 => x"06",
          2931 => x"76",
          2932 => x"3f",
          2933 => x"86",
          2934 => x"f6",
          2935 => x"02",
          2936 => x"05",
          2937 => x"05",
          2938 => x"82",
          2939 => x"70",
          2940 => x"84",
          2941 => x"51",
          2942 => x"58",
          2943 => x"2e",
          2944 => x"51",
          2945 => x"82",
          2946 => x"70",
          2947 => x"84",
          2948 => x"1a",
          2949 => x"51",
          2950 => x"88",
          2951 => x"ec",
          2952 => x"82",
          2953 => x"70",
          2954 => x"84",
          2955 => x"51",
          2956 => x"80",
          2957 => x"75",
          2958 => x"74",
          2959 => x"da",
          2960 => x"c4",
          2961 => x"55",
          2962 => x"c4",
          2963 => x"ff",
          2964 => x"75",
          2965 => x"80",
          2966 => x"c4",
          2967 => x"2e",
          2968 => x"85",
          2969 => x"75",
          2970 => x"38",
          2971 => x"33",
          2972 => x"38",
          2973 => x"05",
          2974 => x"78",
          2975 => x"80",
          2976 => x"82",
          2977 => x"52",
          2978 => x"8a",
          2979 => x"85",
          2980 => x"80",
          2981 => x"8c",
          2982 => x"fd",
          2983 => x"84",
          2984 => x"54",
          2985 => x"71",
          2986 => x"38",
          2987 => x"dd",
          2988 => x"0c",
          2989 => x"14",
          2990 => x"80",
          2991 => x"80",
          2992 => x"c4",
          2993 => x"c0",
          2994 => x"80",
          2995 => x"71",
          2996 => x"dc",
          2997 => x"c0",
          2998 => x"b1",
          2999 => x"82",
          3000 => x"85",
          3001 => x"dc",
          3002 => x"57",
          3003 => x"85",
          3004 => x"80",
          3005 => x"82",
          3006 => x"80",
          3007 => x"85",
          3008 => x"80",
          3009 => x"3d",
          3010 => x"81",
          3011 => x"82",
          3012 => x"80",
          3013 => x"75",
          3014 => x"9e",
          3015 => x"ec",
          3016 => x"0b",
          3017 => x"08",
          3018 => x"82",
          3019 => x"ff",
          3020 => x"55",
          3021 => x"34",
          3022 => x"52",
          3023 => x"fd",
          3024 => x"f6",
          3025 => x"ff",
          3026 => x"06",
          3027 => x"a6",
          3028 => x"d9",
          3029 => x"3d",
          3030 => x"08",
          3031 => x"70",
          3032 => x"52",
          3033 => x"08",
          3034 => x"d2",
          3035 => x"ec",
          3036 => x"38",
          3037 => x"85",
          3038 => x"55",
          3039 => x"8b",
          3040 => x"56",
          3041 => x"3f",
          3042 => x"08",
          3043 => x"38",
          3044 => x"b4",
          3045 => x"85",
          3046 => x"18",
          3047 => x"0b",
          3048 => x"08",
          3049 => x"82",
          3050 => x"ff",
          3051 => x"55",
          3052 => x"34",
          3053 => x"09",
          3054 => x"72",
          3055 => x"51",
          3056 => x"77",
          3057 => x"73",
          3058 => x"82",
          3059 => x"8c",
          3060 => x"51",
          3061 => x"3f",
          3062 => x"08",
          3063 => x"38",
          3064 => x"51",
          3065 => x"78",
          3066 => x"81",
          3067 => x"75",
          3068 => x"ff",
          3069 => x"79",
          3070 => x"be",
          3071 => x"08",
          3072 => x"ec",
          3073 => x"80",
          3074 => x"85",
          3075 => x"3d",
          3076 => x"3d",
          3077 => x"71",
          3078 => x"33",
          3079 => x"58",
          3080 => x"09",
          3081 => x"38",
          3082 => x"05",
          3083 => x"27",
          3084 => x"17",
          3085 => x"71",
          3086 => x"55",
          3087 => x"09",
          3088 => x"38",
          3089 => x"ea",
          3090 => x"74",
          3091 => x"85",
          3092 => x"08",
          3093 => x"ff",
          3094 => x"82",
          3095 => x"53",
          3096 => x"08",
          3097 => x"df",
          3098 => x"ec",
          3099 => x"38",
          3100 => x"54",
          3101 => x"88",
          3102 => x"2e",
          3103 => x"39",
          3104 => x"be",
          3105 => x"5a",
          3106 => x"11",
          3107 => x"51",
          3108 => x"82",
          3109 => x"80",
          3110 => x"ff",
          3111 => x"52",
          3112 => x"af",
          3113 => x"ec",
          3114 => x"06",
          3115 => x"2e",
          3116 => x"15",
          3117 => x"06",
          3118 => x"75",
          3119 => x"38",
          3120 => x"82",
          3121 => x"8c",
          3122 => x"d3",
          3123 => x"3d",
          3124 => x"08",
          3125 => x"59",
          3126 => x"0b",
          3127 => x"82",
          3128 => x"82",
          3129 => x"55",
          3130 => x"ca",
          3131 => x"85",
          3132 => x"55",
          3133 => x"81",
          3134 => x"2e",
          3135 => x"81",
          3136 => x"55",
          3137 => x"2e",
          3138 => x"a8",
          3139 => x"3f",
          3140 => x"08",
          3141 => x"0c",
          3142 => x"08",
          3143 => x"91",
          3144 => x"76",
          3145 => x"ec",
          3146 => x"c8",
          3147 => x"85",
          3148 => x"2e",
          3149 => x"fe",
          3150 => x"a0",
          3151 => x"39",
          3152 => x"08",
          3153 => x"c0",
          3154 => x"f8",
          3155 => x"70",
          3156 => x"82",
          3157 => x"85",
          3158 => x"82",
          3159 => x"74",
          3160 => x"06",
          3161 => x"82",
          3162 => x"51",
          3163 => x"3f",
          3164 => x"08",
          3165 => x"82",
          3166 => x"25",
          3167 => x"85",
          3168 => x"05",
          3169 => x"55",
          3170 => x"80",
          3171 => x"ff",
          3172 => x"51",
          3173 => x"81",
          3174 => x"ff",
          3175 => x"93",
          3176 => x"38",
          3177 => x"ff",
          3178 => x"06",
          3179 => x"86",
          3180 => x"85",
          3181 => x"8c",
          3182 => x"c0",
          3183 => x"84",
          3184 => x"3f",
          3185 => x"e0",
          3186 => x"85",
          3187 => x"2b",
          3188 => x"51",
          3189 => x"2e",
          3190 => x"81",
          3191 => x"9d",
          3192 => x"98",
          3193 => x"2c",
          3194 => x"33",
          3195 => x"70",
          3196 => x"98",
          3197 => x"82",
          3198 => x"f4",
          3199 => x"70",
          3200 => x"51",
          3201 => x"51",
          3202 => x"81",
          3203 => x"2e",
          3204 => x"77",
          3205 => x"38",
          3206 => x"98",
          3207 => x"2c",
          3208 => x"80",
          3209 => x"cb",
          3210 => x"74",
          3211 => x"f6",
          3212 => x"85",
          3213 => x"ff",
          3214 => x"80",
          3215 => x"74",
          3216 => x"34",
          3217 => x"39",
          3218 => x"98",
          3219 => x"2c",
          3220 => x"06",
          3221 => x"54",
          3222 => x"97",
          3223 => x"74",
          3224 => x"f5",
          3225 => x"85",
          3226 => x"ff",
          3227 => x"cf",
          3228 => x"80",
          3229 => x"2e",
          3230 => x"81",
          3231 => x"82",
          3232 => x"73",
          3233 => x"98",
          3234 => x"80",
          3235 => x"2b",
          3236 => x"70",
          3237 => x"82",
          3238 => x"f8",
          3239 => x"52",
          3240 => x"58",
          3241 => x"77",
          3242 => x"06",
          3243 => x"81",
          3244 => x"08",
          3245 => x"0b",
          3246 => x"34",
          3247 => x"9d",
          3248 => x"39",
          3249 => x"84",
          3250 => x"9d",
          3251 => x"af",
          3252 => x"7d",
          3253 => x"73",
          3254 => x"e8",
          3255 => x"2b",
          3256 => x"f0",
          3257 => x"82",
          3258 => x"56",
          3259 => x"fd",
          3260 => x"9d",
          3261 => x"75",
          3262 => x"38",
          3263 => x"70",
          3264 => x"55",
          3265 => x"9e",
          3266 => x"54",
          3267 => x"15",
          3268 => x"70",
          3269 => x"98",
          3270 => x"8c",
          3271 => x"56",
          3272 => x"25",
          3273 => x"9d",
          3274 => x"11",
          3275 => x"82",
          3276 => x"73",
          3277 => x"3d",
          3278 => x"82",
          3279 => x"54",
          3280 => x"89",
          3281 => x"54",
          3282 => x"88",
          3283 => x"8c",
          3284 => x"70",
          3285 => x"98",
          3286 => x"88",
          3287 => x"56",
          3288 => x"25",
          3289 => x"1a",
          3290 => x"54",
          3291 => x"81",
          3292 => x"2b",
          3293 => x"82",
          3294 => x"5a",
          3295 => x"76",
          3296 => x"38",
          3297 => x"33",
          3298 => x"70",
          3299 => x"9d",
          3300 => x"51",
          3301 => x"76",
          3302 => x"38",
          3303 => x"ef",
          3304 => x"70",
          3305 => x"98",
          3306 => x"88",
          3307 => x"56",
          3308 => x"24",
          3309 => x"8c",
          3310 => x"34",
          3311 => x"1b",
          3312 => x"8c",
          3313 => x"81",
          3314 => x"f3",
          3315 => x"d9",
          3316 => x"8c",
          3317 => x"ff",
          3318 => x"73",
          3319 => x"e4",
          3320 => x"88",
          3321 => x"54",
          3322 => x"88",
          3323 => x"54",
          3324 => x"8c",
          3325 => x"e6",
          3326 => x"9d",
          3327 => x"98",
          3328 => x"2c",
          3329 => x"33",
          3330 => x"57",
          3331 => x"a4",
          3332 => x"54",
          3333 => x"74",
          3334 => x"51",
          3335 => x"81",
          3336 => x"2b",
          3337 => x"82",
          3338 => x"59",
          3339 => x"75",
          3340 => x"38",
          3341 => x"d7",
          3342 => x"8c",
          3343 => x"2b",
          3344 => x"82",
          3345 => x"57",
          3346 => x"74",
          3347 => x"f4",
          3348 => x"e5",
          3349 => x"15",
          3350 => x"70",
          3351 => x"9d",
          3352 => x"51",
          3353 => x"75",
          3354 => x"fa",
          3355 => x"9d",
          3356 => x"05",
          3357 => x"34",
          3358 => x"93",
          3359 => x"88",
          3360 => x"f7",
          3361 => x"85",
          3362 => x"ff",
          3363 => x"96",
          3364 => x"88",
          3365 => x"80",
          3366 => x"81",
          3367 => x"79",
          3368 => x"3f",
          3369 => x"7a",
          3370 => x"82",
          3371 => x"80",
          3372 => x"88",
          3373 => x"85",
          3374 => x"3d",
          3375 => x"9d",
          3376 => x"73",
          3377 => x"fc",
          3378 => x"e4",
          3379 => x"9d",
          3380 => x"05",
          3381 => x"9d",
          3382 => x"81",
          3383 => x"e3",
          3384 => x"8c",
          3385 => x"88",
          3386 => x"73",
          3387 => x"d4",
          3388 => x"54",
          3389 => x"88",
          3390 => x"2b",
          3391 => x"75",
          3392 => x"56",
          3393 => x"74",
          3394 => x"74",
          3395 => x"14",
          3396 => x"73",
          3397 => x"f7",
          3398 => x"70",
          3399 => x"98",
          3400 => x"88",
          3401 => x"56",
          3402 => x"24",
          3403 => x"51",
          3404 => x"82",
          3405 => x"70",
          3406 => x"98",
          3407 => x"88",
          3408 => x"56",
          3409 => x"24",
          3410 => x"88",
          3411 => x"3f",
          3412 => x"98",
          3413 => x"2c",
          3414 => x"33",
          3415 => x"54",
          3416 => x"e7",
          3417 => x"39",
          3418 => x"33",
          3419 => x"06",
          3420 => x"33",
          3421 => x"74",
          3422 => x"c8",
          3423 => x"54",
          3424 => x"8c",
          3425 => x"70",
          3426 => x"e3",
          3427 => x"9d",
          3428 => x"81",
          3429 => x"9d",
          3430 => x"56",
          3431 => x"26",
          3432 => x"a0",
          3433 => x"8c",
          3434 => x"81",
          3435 => x"ef",
          3436 => x"0b",
          3437 => x"34",
          3438 => x"9d",
          3439 => x"84",
          3440 => x"38",
          3441 => x"08",
          3442 => x"2e",
          3443 => x"51",
          3444 => x"3f",
          3445 => x"08",
          3446 => x"34",
          3447 => x"08",
          3448 => x"81",
          3449 => x"52",
          3450 => x"a9",
          3451 => x"5b",
          3452 => x"7a",
          3453 => x"84",
          3454 => x"11",
          3455 => x"54",
          3456 => x"a7",
          3457 => x"ff",
          3458 => x"82",
          3459 => x"82",
          3460 => x"82",
          3461 => x"81",
          3462 => x"05",
          3463 => x"79",
          3464 => x"f6",
          3465 => x"54",
          3466 => x"73",
          3467 => x"80",
          3468 => x"38",
          3469 => x"a7",
          3470 => x"39",
          3471 => x"09",
          3472 => x"38",
          3473 => x"08",
          3474 => x"2e",
          3475 => x"51",
          3476 => x"3f",
          3477 => x"08",
          3478 => x"34",
          3479 => x"08",
          3480 => x"81",
          3481 => x"52",
          3482 => x"a8",
          3483 => x"c2",
          3484 => x"2b",
          3485 => x"11",
          3486 => x"74",
          3487 => x"38",
          3488 => x"a6",
          3489 => x"85",
          3490 => x"9d",
          3491 => x"85",
          3492 => x"ff",
          3493 => x"53",
          3494 => x"51",
          3495 => x"3f",
          3496 => x"73",
          3497 => x"5b",
          3498 => x"82",
          3499 => x"74",
          3500 => x"9d",
          3501 => x"9d",
          3502 => x"79",
          3503 => x"3f",
          3504 => x"82",
          3505 => x"70",
          3506 => x"82",
          3507 => x"59",
          3508 => x"77",
          3509 => x"38",
          3510 => x"73",
          3511 => x"34",
          3512 => x"33",
          3513 => x"a7",
          3514 => x"39",
          3515 => x"33",
          3516 => x"2e",
          3517 => x"88",
          3518 => x"3f",
          3519 => x"33",
          3520 => x"73",
          3521 => x"34",
          3522 => x"f9",
          3523 => x"df",
          3524 => x"85",
          3525 => x"80",
          3526 => x"e0",
          3527 => x"53",
          3528 => x"df",
          3529 => x"aa",
          3530 => x"85",
          3531 => x"80",
          3532 => x"34",
          3533 => x"81",
          3534 => x"85",
          3535 => x"77",
          3536 => x"76",
          3537 => x"82",
          3538 => x"54",
          3539 => x"34",
          3540 => x"34",
          3541 => x"08",
          3542 => x"22",
          3543 => x"80",
          3544 => x"83",
          3545 => x"70",
          3546 => x"51",
          3547 => x"88",
          3548 => x"89",
          3549 => x"85",
          3550 => x"83",
          3551 => x"e4",
          3552 => x"05",
          3553 => x"77",
          3554 => x"76",
          3555 => x"89",
          3556 => x"ff",
          3557 => x"52",
          3558 => x"72",
          3559 => x"fb",
          3560 => x"82",
          3561 => x"ff",
          3562 => x"51",
          3563 => x"85",
          3564 => x"3d",
          3565 => x"3d",
          3566 => x"05",
          3567 => x"05",
          3568 => x"71",
          3569 => x"e4",
          3570 => x"2b",
          3571 => x"83",
          3572 => x"70",
          3573 => x"33",
          3574 => x"07",
          3575 => x"ae",
          3576 => x"81",
          3577 => x"07",
          3578 => x"53",
          3579 => x"54",
          3580 => x"53",
          3581 => x"77",
          3582 => x"18",
          3583 => x"e4",
          3584 => x"88",
          3585 => x"70",
          3586 => x"74",
          3587 => x"82",
          3588 => x"70",
          3589 => x"81",
          3590 => x"88",
          3591 => x"83",
          3592 => x"f8",
          3593 => x"56",
          3594 => x"73",
          3595 => x"06",
          3596 => x"54",
          3597 => x"82",
          3598 => x"81",
          3599 => x"72",
          3600 => x"82",
          3601 => x"16",
          3602 => x"34",
          3603 => x"34",
          3604 => x"04",
          3605 => x"82",
          3606 => x"02",
          3607 => x"05",
          3608 => x"2b",
          3609 => x"11",
          3610 => x"33",
          3611 => x"71",
          3612 => x"58",
          3613 => x"55",
          3614 => x"84",
          3615 => x"13",
          3616 => x"2b",
          3617 => x"2a",
          3618 => x"52",
          3619 => x"34",
          3620 => x"34",
          3621 => x"08",
          3622 => x"11",
          3623 => x"33",
          3624 => x"71",
          3625 => x"56",
          3626 => x"72",
          3627 => x"33",
          3628 => x"71",
          3629 => x"70",
          3630 => x"56",
          3631 => x"86",
          3632 => x"87",
          3633 => x"85",
          3634 => x"70",
          3635 => x"33",
          3636 => x"07",
          3637 => x"ff",
          3638 => x"2a",
          3639 => x"53",
          3640 => x"34",
          3641 => x"34",
          3642 => x"04",
          3643 => x"02",
          3644 => x"82",
          3645 => x"71",
          3646 => x"11",
          3647 => x"12",
          3648 => x"2b",
          3649 => x"2b",
          3650 => x"55",
          3651 => x"70",
          3652 => x"33",
          3653 => x"71",
          3654 => x"53",
          3655 => x"55",
          3656 => x"80",
          3657 => x"51",
          3658 => x"82",
          3659 => x"70",
          3660 => x"81",
          3661 => x"8b",
          3662 => x"2b",
          3663 => x"70",
          3664 => x"33",
          3665 => x"07",
          3666 => x"8f",
          3667 => x"51",
          3668 => x"53",
          3669 => x"72",
          3670 => x"2a",
          3671 => x"82",
          3672 => x"83",
          3673 => x"85",
          3674 => x"17",
          3675 => x"12",
          3676 => x"2b",
          3677 => x"07",
          3678 => x"55",
          3679 => x"33",
          3680 => x"71",
          3681 => x"70",
          3682 => x"06",
          3683 => x"57",
          3684 => x"52",
          3685 => x"71",
          3686 => x"89",
          3687 => x"fb",
          3688 => x"85",
          3689 => x"84",
          3690 => x"22",
          3691 => x"72",
          3692 => x"33",
          3693 => x"71",
          3694 => x"83",
          3695 => x"5b",
          3696 => x"52",
          3697 => x"33",
          3698 => x"71",
          3699 => x"02",
          3700 => x"05",
          3701 => x"70",
          3702 => x"51",
          3703 => x"71",
          3704 => x"81",
          3705 => x"85",
          3706 => x"15",
          3707 => x"12",
          3708 => x"2b",
          3709 => x"07",
          3710 => x"52",
          3711 => x"12",
          3712 => x"33",
          3713 => x"07",
          3714 => x"54",
          3715 => x"70",
          3716 => x"72",
          3717 => x"82",
          3718 => x"14",
          3719 => x"83",
          3720 => x"88",
          3721 => x"85",
          3722 => x"54",
          3723 => x"04",
          3724 => x"7b",
          3725 => x"08",
          3726 => x"70",
          3727 => x"06",
          3728 => x"53",
          3729 => x"82",
          3730 => x"76",
          3731 => x"11",
          3732 => x"83",
          3733 => x"8b",
          3734 => x"2b",
          3735 => x"70",
          3736 => x"33",
          3737 => x"71",
          3738 => x"53",
          3739 => x"53",
          3740 => x"59",
          3741 => x"25",
          3742 => x"80",
          3743 => x"51",
          3744 => x"81",
          3745 => x"14",
          3746 => x"33",
          3747 => x"71",
          3748 => x"76",
          3749 => x"2a",
          3750 => x"58",
          3751 => x"14",
          3752 => x"ff",
          3753 => x"87",
          3754 => x"85",
          3755 => x"19",
          3756 => x"85",
          3757 => x"88",
          3758 => x"88",
          3759 => x"5b",
          3760 => x"84",
          3761 => x"85",
          3762 => x"85",
          3763 => x"53",
          3764 => x"14",
          3765 => x"87",
          3766 => x"85",
          3767 => x"76",
          3768 => x"75",
          3769 => x"82",
          3770 => x"18",
          3771 => x"12",
          3772 => x"2b",
          3773 => x"80",
          3774 => x"88",
          3775 => x"55",
          3776 => x"74",
          3777 => x"15",
          3778 => x"0d",
          3779 => x"0d",
          3780 => x"85",
          3781 => x"38",
          3782 => x"71",
          3783 => x"38",
          3784 => x"8c",
          3785 => x"0d",
          3786 => x"0d",
          3787 => x"58",
          3788 => x"82",
          3789 => x"83",
          3790 => x"82",
          3791 => x"84",
          3792 => x"12",
          3793 => x"2b",
          3794 => x"59",
          3795 => x"81",
          3796 => x"75",
          3797 => x"cc",
          3798 => x"2b",
          3799 => x"33",
          3800 => x"71",
          3801 => x"70",
          3802 => x"06",
          3803 => x"83",
          3804 => x"70",
          3805 => x"53",
          3806 => x"55",
          3807 => x"8a",
          3808 => x"2e",
          3809 => x"78",
          3810 => x"15",
          3811 => x"33",
          3812 => x"07",
          3813 => x"c1",
          3814 => x"ff",
          3815 => x"38",
          3816 => x"56",
          3817 => x"2b",
          3818 => x"08",
          3819 => x"81",
          3820 => x"88",
          3821 => x"81",
          3822 => x"51",
          3823 => x"5c",
          3824 => x"2e",
          3825 => x"55",
          3826 => x"78",
          3827 => x"38",
          3828 => x"80",
          3829 => x"38",
          3830 => x"09",
          3831 => x"38",
          3832 => x"f0",
          3833 => x"39",
          3834 => x"53",
          3835 => x"51",
          3836 => x"82",
          3837 => x"70",
          3838 => x"33",
          3839 => x"71",
          3840 => x"83",
          3841 => x"5a",
          3842 => x"05",
          3843 => x"83",
          3844 => x"70",
          3845 => x"59",
          3846 => x"84",
          3847 => x"81",
          3848 => x"76",
          3849 => x"82",
          3850 => x"75",
          3851 => x"11",
          3852 => x"11",
          3853 => x"33",
          3854 => x"07",
          3855 => x"53",
          3856 => x"5a",
          3857 => x"86",
          3858 => x"87",
          3859 => x"85",
          3860 => x"1c",
          3861 => x"85",
          3862 => x"8b",
          3863 => x"2b",
          3864 => x"5a",
          3865 => x"54",
          3866 => x"34",
          3867 => x"34",
          3868 => x"08",
          3869 => x"1d",
          3870 => x"85",
          3871 => x"88",
          3872 => x"88",
          3873 => x"5f",
          3874 => x"73",
          3875 => x"75",
          3876 => x"82",
          3877 => x"1b",
          3878 => x"73",
          3879 => x"0c",
          3880 => x"04",
          3881 => x"74",
          3882 => x"e4",
          3883 => x"f4",
          3884 => x"53",
          3885 => x"8b",
          3886 => x"fc",
          3887 => x"85",
          3888 => x"72",
          3889 => x"0c",
          3890 => x"04",
          3891 => x"02",
          3892 => x"51",
          3893 => x"72",
          3894 => x"82",
          3895 => x"33",
          3896 => x"85",
          3897 => x"3d",
          3898 => x"3d",
          3899 => x"05",
          3900 => x"05",
          3901 => x"56",
          3902 => x"72",
          3903 => x"e0",
          3904 => x"2b",
          3905 => x"8c",
          3906 => x"88",
          3907 => x"2e",
          3908 => x"88",
          3909 => x"0c",
          3910 => x"8c",
          3911 => x"71",
          3912 => x"87",
          3913 => x"0c",
          3914 => x"08",
          3915 => x"51",
          3916 => x"2e",
          3917 => x"c0",
          3918 => x"51",
          3919 => x"71",
          3920 => x"80",
          3921 => x"92",
          3922 => x"98",
          3923 => x"70",
          3924 => x"38",
          3925 => x"e8",
          3926 => x"85",
          3927 => x"51",
          3928 => x"ec",
          3929 => x"0d",
          3930 => x"0d",
          3931 => x"02",
          3932 => x"05",
          3933 => x"58",
          3934 => x"52",
          3935 => x"3f",
          3936 => x"08",
          3937 => x"54",
          3938 => x"be",
          3939 => x"75",
          3940 => x"c0",
          3941 => x"87",
          3942 => x"12",
          3943 => x"84",
          3944 => x"40",
          3945 => x"85",
          3946 => x"98",
          3947 => x"7d",
          3948 => x"0c",
          3949 => x"85",
          3950 => x"06",
          3951 => x"71",
          3952 => x"38",
          3953 => x"71",
          3954 => x"05",
          3955 => x"19",
          3956 => x"a2",
          3957 => x"71",
          3958 => x"38",
          3959 => x"83",
          3960 => x"38",
          3961 => x"8a",
          3962 => x"98",
          3963 => x"71",
          3964 => x"c0",
          3965 => x"52",
          3966 => x"87",
          3967 => x"80",
          3968 => x"81",
          3969 => x"c0",
          3970 => x"53",
          3971 => x"82",
          3972 => x"71",
          3973 => x"1a",
          3974 => x"84",
          3975 => x"19",
          3976 => x"06",
          3977 => x"79",
          3978 => x"38",
          3979 => x"80",
          3980 => x"87",
          3981 => x"26",
          3982 => x"73",
          3983 => x"06",
          3984 => x"2e",
          3985 => x"52",
          3986 => x"82",
          3987 => x"8f",
          3988 => x"f3",
          3989 => x"62",
          3990 => x"05",
          3991 => x"57",
          3992 => x"83",
          3993 => x"52",
          3994 => x"3f",
          3995 => x"08",
          3996 => x"54",
          3997 => x"2e",
          3998 => x"81",
          3999 => x"74",
          4000 => x"c0",
          4001 => x"87",
          4002 => x"12",
          4003 => x"84",
          4004 => x"5f",
          4005 => x"0b",
          4006 => x"8c",
          4007 => x"0c",
          4008 => x"80",
          4009 => x"70",
          4010 => x"81",
          4011 => x"54",
          4012 => x"8c",
          4013 => x"81",
          4014 => x"7c",
          4015 => x"58",
          4016 => x"70",
          4017 => x"52",
          4018 => x"8a",
          4019 => x"98",
          4020 => x"71",
          4021 => x"c0",
          4022 => x"52",
          4023 => x"87",
          4024 => x"80",
          4025 => x"81",
          4026 => x"c0",
          4027 => x"53",
          4028 => x"82",
          4029 => x"71",
          4030 => x"19",
          4031 => x"81",
          4032 => x"ff",
          4033 => x"19",
          4034 => x"78",
          4035 => x"38",
          4036 => x"80",
          4037 => x"87",
          4038 => x"26",
          4039 => x"73",
          4040 => x"06",
          4041 => x"2e",
          4042 => x"52",
          4043 => x"82",
          4044 => x"8f",
          4045 => x"fa",
          4046 => x"02",
          4047 => x"05",
          4048 => x"05",
          4049 => x"71",
          4050 => x"57",
          4051 => x"82",
          4052 => x"81",
          4053 => x"54",
          4054 => x"38",
          4055 => x"c0",
          4056 => x"81",
          4057 => x"2e",
          4058 => x"71",
          4059 => x"38",
          4060 => x"87",
          4061 => x"11",
          4062 => x"80",
          4063 => x"80",
          4064 => x"83",
          4065 => x"38",
          4066 => x"72",
          4067 => x"2a",
          4068 => x"51",
          4069 => x"80",
          4070 => x"87",
          4071 => x"08",
          4072 => x"38",
          4073 => x"8c",
          4074 => x"96",
          4075 => x"0c",
          4076 => x"8c",
          4077 => x"08",
          4078 => x"51",
          4079 => x"38",
          4080 => x"56",
          4081 => x"80",
          4082 => x"85",
          4083 => x"77",
          4084 => x"83",
          4085 => x"75",
          4086 => x"85",
          4087 => x"3d",
          4088 => x"3d",
          4089 => x"11",
          4090 => x"71",
          4091 => x"82",
          4092 => x"53",
          4093 => x"0d",
          4094 => x"0d",
          4095 => x"33",
          4096 => x"71",
          4097 => x"88",
          4098 => x"14",
          4099 => x"07",
          4100 => x"33",
          4101 => x"85",
          4102 => x"53",
          4103 => x"52",
          4104 => x"04",
          4105 => x"73",
          4106 => x"92",
          4107 => x"52",
          4108 => x"81",
          4109 => x"70",
          4110 => x"70",
          4111 => x"3d",
          4112 => x"3d",
          4113 => x"52",
          4114 => x"70",
          4115 => x"34",
          4116 => x"51",
          4117 => x"81",
          4118 => x"70",
          4119 => x"70",
          4120 => x"05",
          4121 => x"88",
          4122 => x"72",
          4123 => x"0d",
          4124 => x"0d",
          4125 => x"54",
          4126 => x"80",
          4127 => x"71",
          4128 => x"53",
          4129 => x"81",
          4130 => x"ff",
          4131 => x"39",
          4132 => x"04",
          4133 => x"75",
          4134 => x"52",
          4135 => x"70",
          4136 => x"34",
          4137 => x"70",
          4138 => x"3d",
          4139 => x"3d",
          4140 => x"79",
          4141 => x"74",
          4142 => x"56",
          4143 => x"81",
          4144 => x"71",
          4145 => x"16",
          4146 => x"52",
          4147 => x"86",
          4148 => x"2e",
          4149 => x"82",
          4150 => x"86",
          4151 => x"fe",
          4152 => x"76",
          4153 => x"39",
          4154 => x"8a",
          4155 => x"51",
          4156 => x"71",
          4157 => x"33",
          4158 => x"0c",
          4159 => x"04",
          4160 => x"85",
          4161 => x"80",
          4162 => x"ec",
          4163 => x"3d",
          4164 => x"80",
          4165 => x"33",
          4166 => x"7a",
          4167 => x"38",
          4168 => x"16",
          4169 => x"16",
          4170 => x"17",
          4171 => x"fa",
          4172 => x"85",
          4173 => x"2e",
          4174 => x"b7",
          4175 => x"ec",
          4176 => x"34",
          4177 => x"70",
          4178 => x"31",
          4179 => x"59",
          4180 => x"77",
          4181 => x"82",
          4182 => x"74",
          4183 => x"81",
          4184 => x"81",
          4185 => x"53",
          4186 => x"16",
          4187 => x"e3",
          4188 => x"81",
          4189 => x"85",
          4190 => x"3d",
          4191 => x"3d",
          4192 => x"56",
          4193 => x"74",
          4194 => x"2e",
          4195 => x"51",
          4196 => x"82",
          4197 => x"57",
          4198 => x"08",
          4199 => x"54",
          4200 => x"16",
          4201 => x"33",
          4202 => x"3f",
          4203 => x"08",
          4204 => x"38",
          4205 => x"57",
          4206 => x"0c",
          4207 => x"ec",
          4208 => x"0d",
          4209 => x"0d",
          4210 => x"57",
          4211 => x"82",
          4212 => x"58",
          4213 => x"08",
          4214 => x"76",
          4215 => x"83",
          4216 => x"06",
          4217 => x"84",
          4218 => x"78",
          4219 => x"81",
          4220 => x"38",
          4221 => x"82",
          4222 => x"52",
          4223 => x"52",
          4224 => x"3f",
          4225 => x"52",
          4226 => x"51",
          4227 => x"84",
          4228 => x"d2",
          4229 => x"fc",
          4230 => x"8a",
          4231 => x"52",
          4232 => x"51",
          4233 => x"90",
          4234 => x"84",
          4235 => x"fc",
          4236 => x"17",
          4237 => x"a0",
          4238 => x"86",
          4239 => x"08",
          4240 => x"b0",
          4241 => x"55",
          4242 => x"81",
          4243 => x"f8",
          4244 => x"84",
          4245 => x"53",
          4246 => x"17",
          4247 => x"d7",
          4248 => x"ec",
          4249 => x"83",
          4250 => x"77",
          4251 => x"0c",
          4252 => x"04",
          4253 => x"77",
          4254 => x"12",
          4255 => x"55",
          4256 => x"56",
          4257 => x"94",
          4258 => x"22",
          4259 => x"ff",
          4260 => x"ac",
          4261 => x"85",
          4262 => x"56",
          4263 => x"ec",
          4264 => x"0d",
          4265 => x"0d",
          4266 => x"08",
          4267 => x"81",
          4268 => x"df",
          4269 => x"15",
          4270 => x"d7",
          4271 => x"33",
          4272 => x"82",
          4273 => x"38",
          4274 => x"89",
          4275 => x"2e",
          4276 => x"bf",
          4277 => x"2e",
          4278 => x"81",
          4279 => x"81",
          4280 => x"89",
          4281 => x"08",
          4282 => x"52",
          4283 => x"3f",
          4284 => x"08",
          4285 => x"74",
          4286 => x"14",
          4287 => x"81",
          4288 => x"2a",
          4289 => x"05",
          4290 => x"57",
          4291 => x"ee",
          4292 => x"ec",
          4293 => x"38",
          4294 => x"06",
          4295 => x"33",
          4296 => x"78",
          4297 => x"06",
          4298 => x"5c",
          4299 => x"53",
          4300 => x"38",
          4301 => x"06",
          4302 => x"39",
          4303 => x"a4",
          4304 => x"52",
          4305 => x"b6",
          4306 => x"ec",
          4307 => x"38",
          4308 => x"fe",
          4309 => x"b4",
          4310 => x"86",
          4311 => x"ec",
          4312 => x"ff",
          4313 => x"39",
          4314 => x"a4",
          4315 => x"52",
          4316 => x"8a",
          4317 => x"ec",
          4318 => x"76",
          4319 => x"fc",
          4320 => x"b4",
          4321 => x"f1",
          4322 => x"ec",
          4323 => x"06",
          4324 => x"81",
          4325 => x"85",
          4326 => x"3d",
          4327 => x"3d",
          4328 => x"7e",
          4329 => x"82",
          4330 => x"27",
          4331 => x"76",
          4332 => x"27",
          4333 => x"75",
          4334 => x"79",
          4335 => x"38",
          4336 => x"89",
          4337 => x"2e",
          4338 => x"80",
          4339 => x"2e",
          4340 => x"81",
          4341 => x"81",
          4342 => x"89",
          4343 => x"08",
          4344 => x"52",
          4345 => x"3f",
          4346 => x"08",
          4347 => x"ec",
          4348 => x"38",
          4349 => x"06",
          4350 => x"81",
          4351 => x"06",
          4352 => x"77",
          4353 => x"2e",
          4354 => x"84",
          4355 => x"06",
          4356 => x"06",
          4357 => x"53",
          4358 => x"81",
          4359 => x"34",
          4360 => x"a4",
          4361 => x"52",
          4362 => x"d2",
          4363 => x"ec",
          4364 => x"85",
          4365 => x"94",
          4366 => x"ff",
          4367 => x"05",
          4368 => x"54",
          4369 => x"38",
          4370 => x"74",
          4371 => x"06",
          4372 => x"07",
          4373 => x"74",
          4374 => x"39",
          4375 => x"a4",
          4376 => x"52",
          4377 => x"96",
          4378 => x"ec",
          4379 => x"85",
          4380 => x"d8",
          4381 => x"ff",
          4382 => x"76",
          4383 => x"06",
          4384 => x"05",
          4385 => x"3f",
          4386 => x"87",
          4387 => x"08",
          4388 => x"51",
          4389 => x"82",
          4390 => x"59",
          4391 => x"08",
          4392 => x"f0",
          4393 => x"82",
          4394 => x"06",
          4395 => x"05",
          4396 => x"54",
          4397 => x"3f",
          4398 => x"08",
          4399 => x"74",
          4400 => x"51",
          4401 => x"81",
          4402 => x"34",
          4403 => x"ec",
          4404 => x"0d",
          4405 => x"0d",
          4406 => x"72",
          4407 => x"56",
          4408 => x"27",
          4409 => x"98",
          4410 => x"9d",
          4411 => x"2e",
          4412 => x"53",
          4413 => x"51",
          4414 => x"82",
          4415 => x"54",
          4416 => x"08",
          4417 => x"93",
          4418 => x"80",
          4419 => x"54",
          4420 => x"82",
          4421 => x"54",
          4422 => x"74",
          4423 => x"fb",
          4424 => x"85",
          4425 => x"82",
          4426 => x"80",
          4427 => x"38",
          4428 => x"08",
          4429 => x"38",
          4430 => x"08",
          4431 => x"38",
          4432 => x"52",
          4433 => x"d6",
          4434 => x"ec",
          4435 => x"98",
          4436 => x"11",
          4437 => x"57",
          4438 => x"74",
          4439 => x"81",
          4440 => x"0c",
          4441 => x"81",
          4442 => x"84",
          4443 => x"55",
          4444 => x"ff",
          4445 => x"54",
          4446 => x"ec",
          4447 => x"0d",
          4448 => x"0d",
          4449 => x"08",
          4450 => x"79",
          4451 => x"17",
          4452 => x"80",
          4453 => x"98",
          4454 => x"26",
          4455 => x"58",
          4456 => x"52",
          4457 => x"fd",
          4458 => x"74",
          4459 => x"08",
          4460 => x"38",
          4461 => x"08",
          4462 => x"ec",
          4463 => x"82",
          4464 => x"17",
          4465 => x"ec",
          4466 => x"cd",
          4467 => x"90",
          4468 => x"56",
          4469 => x"2e",
          4470 => x"77",
          4471 => x"81",
          4472 => x"38",
          4473 => x"98",
          4474 => x"26",
          4475 => x"56",
          4476 => x"51",
          4477 => x"80",
          4478 => x"ec",
          4479 => x"09",
          4480 => x"38",
          4481 => x"08",
          4482 => x"ec",
          4483 => x"09",
          4484 => x"72",
          4485 => x"70",
          4486 => x"85",
          4487 => x"51",
          4488 => x"73",
          4489 => x"82",
          4490 => x"80",
          4491 => x"8c",
          4492 => x"81",
          4493 => x"38",
          4494 => x"08",
          4495 => x"73",
          4496 => x"75",
          4497 => x"77",
          4498 => x"56",
          4499 => x"76",
          4500 => x"82",
          4501 => x"26",
          4502 => x"75",
          4503 => x"f8",
          4504 => x"85",
          4505 => x"2e",
          4506 => x"59",
          4507 => x"08",
          4508 => x"81",
          4509 => x"82",
          4510 => x"59",
          4511 => x"08",
          4512 => x"81",
          4513 => x"07",
          4514 => x"7c",
          4515 => x"55",
          4516 => x"fa",
          4517 => x"2e",
          4518 => x"ff",
          4519 => x"55",
          4520 => x"ff",
          4521 => x"76",
          4522 => x"3f",
          4523 => x"08",
          4524 => x"08",
          4525 => x"70",
          4526 => x"08",
          4527 => x"51",
          4528 => x"80",
          4529 => x"73",
          4530 => x"38",
          4531 => x"52",
          4532 => x"ca",
          4533 => x"ec",
          4534 => x"a5",
          4535 => x"18",
          4536 => x"08",
          4537 => x"18",
          4538 => x"74",
          4539 => x"38",
          4540 => x"18",
          4541 => x"33",
          4542 => x"73",
          4543 => x"97",
          4544 => x"74",
          4545 => x"38",
          4546 => x"55",
          4547 => x"85",
          4548 => x"85",
          4549 => x"75",
          4550 => x"85",
          4551 => x"3d",
          4552 => x"3d",
          4553 => x"52",
          4554 => x"3f",
          4555 => x"08",
          4556 => x"82",
          4557 => x"80",
          4558 => x"52",
          4559 => x"b4",
          4560 => x"ec",
          4561 => x"ec",
          4562 => x"0c",
          4563 => x"53",
          4564 => x"15",
          4565 => x"f2",
          4566 => x"56",
          4567 => x"16",
          4568 => x"22",
          4569 => x"27",
          4570 => x"54",
          4571 => x"76",
          4572 => x"33",
          4573 => x"3f",
          4574 => x"08",
          4575 => x"38",
          4576 => x"76",
          4577 => x"81",
          4578 => x"07",
          4579 => x"53",
          4580 => x"75",
          4581 => x"0c",
          4582 => x"04",
          4583 => x"7a",
          4584 => x"58",
          4585 => x"f0",
          4586 => x"80",
          4587 => x"9f",
          4588 => x"80",
          4589 => x"90",
          4590 => x"17",
          4591 => x"aa",
          4592 => x"53",
          4593 => x"88",
          4594 => x"08",
          4595 => x"38",
          4596 => x"53",
          4597 => x"17",
          4598 => x"72",
          4599 => x"fe",
          4600 => x"08",
          4601 => x"80",
          4602 => x"16",
          4603 => x"2b",
          4604 => x"75",
          4605 => x"73",
          4606 => x"f5",
          4607 => x"85",
          4608 => x"82",
          4609 => x"ff",
          4610 => x"81",
          4611 => x"ec",
          4612 => x"38",
          4613 => x"82",
          4614 => x"26",
          4615 => x"58",
          4616 => x"73",
          4617 => x"39",
          4618 => x"51",
          4619 => x"82",
          4620 => x"98",
          4621 => x"94",
          4622 => x"17",
          4623 => x"58",
          4624 => x"9a",
          4625 => x"81",
          4626 => x"74",
          4627 => x"98",
          4628 => x"83",
          4629 => x"b4",
          4630 => x"0c",
          4631 => x"82",
          4632 => x"8a",
          4633 => x"f8",
          4634 => x"70",
          4635 => x"08",
          4636 => x"57",
          4637 => x"0a",
          4638 => x"38",
          4639 => x"15",
          4640 => x"08",
          4641 => x"72",
          4642 => x"cb",
          4643 => x"ff",
          4644 => x"81",
          4645 => x"13",
          4646 => x"94",
          4647 => x"74",
          4648 => x"85",
          4649 => x"22",
          4650 => x"73",
          4651 => x"38",
          4652 => x"8a",
          4653 => x"05",
          4654 => x"06",
          4655 => x"8a",
          4656 => x"73",
          4657 => x"3f",
          4658 => x"08",
          4659 => x"81",
          4660 => x"ec",
          4661 => x"ff",
          4662 => x"82",
          4663 => x"ff",
          4664 => x"38",
          4665 => x"82",
          4666 => x"26",
          4667 => x"7b",
          4668 => x"98",
          4669 => x"55",
          4670 => x"94",
          4671 => x"73",
          4672 => x"3f",
          4673 => x"08",
          4674 => x"82",
          4675 => x"80",
          4676 => x"38",
          4677 => x"85",
          4678 => x"2e",
          4679 => x"55",
          4680 => x"08",
          4681 => x"38",
          4682 => x"08",
          4683 => x"fb",
          4684 => x"85",
          4685 => x"38",
          4686 => x"0c",
          4687 => x"51",
          4688 => x"82",
          4689 => x"98",
          4690 => x"90",
          4691 => x"16",
          4692 => x"15",
          4693 => x"74",
          4694 => x"0c",
          4695 => x"04",
          4696 => x"7b",
          4697 => x"5b",
          4698 => x"52",
          4699 => x"ac",
          4700 => x"ec",
          4701 => x"85",
          4702 => x"ec",
          4703 => x"ec",
          4704 => x"17",
          4705 => x"51",
          4706 => x"82",
          4707 => x"54",
          4708 => x"08",
          4709 => x"82",
          4710 => x"9c",
          4711 => x"33",
          4712 => x"72",
          4713 => x"09",
          4714 => x"38",
          4715 => x"85",
          4716 => x"72",
          4717 => x"55",
          4718 => x"53",
          4719 => x"8e",
          4720 => x"56",
          4721 => x"09",
          4722 => x"38",
          4723 => x"85",
          4724 => x"81",
          4725 => x"fd",
          4726 => x"85",
          4727 => x"82",
          4728 => x"80",
          4729 => x"38",
          4730 => x"09",
          4731 => x"38",
          4732 => x"82",
          4733 => x"8b",
          4734 => x"fd",
          4735 => x"9a",
          4736 => x"eb",
          4737 => x"85",
          4738 => x"ff",
          4739 => x"70",
          4740 => x"53",
          4741 => x"09",
          4742 => x"38",
          4743 => x"eb",
          4744 => x"85",
          4745 => x"2b",
          4746 => x"72",
          4747 => x"0c",
          4748 => x"04",
          4749 => x"77",
          4750 => x"ff",
          4751 => x"9a",
          4752 => x"55",
          4753 => x"76",
          4754 => x"53",
          4755 => x"09",
          4756 => x"38",
          4757 => x"52",
          4758 => x"eb",
          4759 => x"3d",
          4760 => x"3d",
          4761 => x"5b",
          4762 => x"08",
          4763 => x"15",
          4764 => x"81",
          4765 => x"15",
          4766 => x"51",
          4767 => x"82",
          4768 => x"58",
          4769 => x"08",
          4770 => x"9c",
          4771 => x"33",
          4772 => x"86",
          4773 => x"80",
          4774 => x"13",
          4775 => x"06",
          4776 => x"06",
          4777 => x"72",
          4778 => x"82",
          4779 => x"53",
          4780 => x"2e",
          4781 => x"53",
          4782 => x"a9",
          4783 => x"74",
          4784 => x"72",
          4785 => x"38",
          4786 => x"99",
          4787 => x"ec",
          4788 => x"06",
          4789 => x"88",
          4790 => x"06",
          4791 => x"54",
          4792 => x"a0",
          4793 => x"74",
          4794 => x"3f",
          4795 => x"08",
          4796 => x"ec",
          4797 => x"98",
          4798 => x"fa",
          4799 => x"80",
          4800 => x"0c",
          4801 => x"ec",
          4802 => x"0d",
          4803 => x"0d",
          4804 => x"57",
          4805 => x"73",
          4806 => x"3f",
          4807 => x"08",
          4808 => x"ec",
          4809 => x"98",
          4810 => x"75",
          4811 => x"3f",
          4812 => x"08",
          4813 => x"ec",
          4814 => x"a0",
          4815 => x"ec",
          4816 => x"14",
          4817 => x"cc",
          4818 => x"a0",
          4819 => x"14",
          4820 => x"9d",
          4821 => x"83",
          4822 => x"82",
          4823 => x"87",
          4824 => x"fd",
          4825 => x"70",
          4826 => x"08",
          4827 => x"55",
          4828 => x"3f",
          4829 => x"08",
          4830 => x"13",
          4831 => x"73",
          4832 => x"83",
          4833 => x"3d",
          4834 => x"3d",
          4835 => x"57",
          4836 => x"89",
          4837 => x"17",
          4838 => x"81",
          4839 => x"70",
          4840 => x"55",
          4841 => x"08",
          4842 => x"81",
          4843 => x"52",
          4844 => x"a8",
          4845 => x"2e",
          4846 => x"84",
          4847 => x"52",
          4848 => x"09",
          4849 => x"38",
          4850 => x"81",
          4851 => x"81",
          4852 => x"73",
          4853 => x"55",
          4854 => x"55",
          4855 => x"c5",
          4856 => x"88",
          4857 => x"0b",
          4858 => x"9c",
          4859 => x"8b",
          4860 => x"17",
          4861 => x"08",
          4862 => x"52",
          4863 => x"82",
          4864 => x"76",
          4865 => x"51",
          4866 => x"82",
          4867 => x"86",
          4868 => x"12",
          4869 => x"3f",
          4870 => x"08",
          4871 => x"88",
          4872 => x"f3",
          4873 => x"70",
          4874 => x"80",
          4875 => x"51",
          4876 => x"af",
          4877 => x"81",
          4878 => x"dc",
          4879 => x"74",
          4880 => x"38",
          4881 => x"88",
          4882 => x"39",
          4883 => x"80",
          4884 => x"56",
          4885 => x"af",
          4886 => x"06",
          4887 => x"56",
          4888 => x"32",
          4889 => x"05",
          4890 => x"78",
          4891 => x"54",
          4892 => x"73",
          4893 => x"60",
          4894 => x"54",
          4895 => x"96",
          4896 => x"0b",
          4897 => x"80",
          4898 => x"f6",
          4899 => x"85",
          4900 => x"85",
          4901 => x"3d",
          4902 => x"5c",
          4903 => x"53",
          4904 => x"51",
          4905 => x"80",
          4906 => x"88",
          4907 => x"5c",
          4908 => x"09",
          4909 => x"d8",
          4910 => x"70",
          4911 => x"71",
          4912 => x"09",
          4913 => x"9f",
          4914 => x"26",
          4915 => x"53",
          4916 => x"73",
          4917 => x"17",
          4918 => x"34",
          4919 => x"d9",
          4920 => x"32",
          4921 => x"05",
          4922 => x"51",
          4923 => x"80",
          4924 => x"38",
          4925 => x"87",
          4926 => x"26",
          4927 => x"77",
          4928 => x"a4",
          4929 => x"27",
          4930 => x"a0",
          4931 => x"39",
          4932 => x"33",
          4933 => x"57",
          4934 => x"27",
          4935 => x"75",
          4936 => x"09",
          4937 => x"80",
          4938 => x"09",
          4939 => x"80",
          4940 => x"25",
          4941 => x"56",
          4942 => x"80",
          4943 => x"84",
          4944 => x"58",
          4945 => x"70",
          4946 => x"55",
          4947 => x"09",
          4948 => x"38",
          4949 => x"80",
          4950 => x"09",
          4951 => x"80",
          4952 => x"51",
          4953 => x"d9",
          4954 => x"39",
          4955 => x"09",
          4956 => x"38",
          4957 => x"7c",
          4958 => x"54",
          4959 => x"a6",
          4960 => x"32",
          4961 => x"05",
          4962 => x"70",
          4963 => x"72",
          4964 => x"9f",
          4965 => x"51",
          4966 => x"74",
          4967 => x"88",
          4968 => x"fe",
          4969 => x"98",
          4970 => x"80",
          4971 => x"75",
          4972 => x"81",
          4973 => x"33",
          4974 => x"51",
          4975 => x"82",
          4976 => x"80",
          4977 => x"78",
          4978 => x"81",
          4979 => x"5a",
          4980 => x"b3",
          4981 => x"ec",
          4982 => x"80",
          4983 => x"1c",
          4984 => x"27",
          4985 => x"79",
          4986 => x"74",
          4987 => x"7a",
          4988 => x"74",
          4989 => x"39",
          4990 => x"fe",
          4991 => x"df",
          4992 => x"ec",
          4993 => x"ff",
          4994 => x"73",
          4995 => x"38",
          4996 => x"81",
          4997 => x"54",
          4998 => x"75",
          4999 => x"17",
          5000 => x"39",
          5001 => x"0c",
          5002 => x"99",
          5003 => x"54",
          5004 => x"2e",
          5005 => x"84",
          5006 => x"34",
          5007 => x"76",
          5008 => x"8b",
          5009 => x"81",
          5010 => x"56",
          5011 => x"80",
          5012 => x"1b",
          5013 => x"08",
          5014 => x"51",
          5015 => x"82",
          5016 => x"56",
          5017 => x"08",
          5018 => x"98",
          5019 => x"76",
          5020 => x"3f",
          5021 => x"08",
          5022 => x"ec",
          5023 => x"38",
          5024 => x"70",
          5025 => x"73",
          5026 => x"be",
          5027 => x"33",
          5028 => x"73",
          5029 => x"8b",
          5030 => x"83",
          5031 => x"06",
          5032 => x"73",
          5033 => x"53",
          5034 => x"51",
          5035 => x"82",
          5036 => x"80",
          5037 => x"75",
          5038 => x"f3",
          5039 => x"9f",
          5040 => x"1c",
          5041 => x"74",
          5042 => x"38",
          5043 => x"09",
          5044 => x"e7",
          5045 => x"2a",
          5046 => x"77",
          5047 => x"51",
          5048 => x"2e",
          5049 => x"81",
          5050 => x"80",
          5051 => x"38",
          5052 => x"ab",
          5053 => x"55",
          5054 => x"75",
          5055 => x"73",
          5056 => x"55",
          5057 => x"82",
          5058 => x"06",
          5059 => x"ab",
          5060 => x"33",
          5061 => x"70",
          5062 => x"55",
          5063 => x"2e",
          5064 => x"1b",
          5065 => x"06",
          5066 => x"52",
          5067 => x"cb",
          5068 => x"ec",
          5069 => x"0c",
          5070 => x"74",
          5071 => x"0c",
          5072 => x"04",
          5073 => x"7c",
          5074 => x"08",
          5075 => x"55",
          5076 => x"59",
          5077 => x"81",
          5078 => x"70",
          5079 => x"33",
          5080 => x"52",
          5081 => x"2e",
          5082 => x"ee",
          5083 => x"2e",
          5084 => x"81",
          5085 => x"33",
          5086 => x"81",
          5087 => x"52",
          5088 => x"26",
          5089 => x"14",
          5090 => x"06",
          5091 => x"52",
          5092 => x"80",
          5093 => x"0b",
          5094 => x"59",
          5095 => x"7a",
          5096 => x"70",
          5097 => x"33",
          5098 => x"05",
          5099 => x"9f",
          5100 => x"53",
          5101 => x"89",
          5102 => x"70",
          5103 => x"54",
          5104 => x"12",
          5105 => x"26",
          5106 => x"12",
          5107 => x"06",
          5108 => x"09",
          5109 => x"9f",
          5110 => x"72",
          5111 => x"81",
          5112 => x"70",
          5113 => x"72",
          5114 => x"74",
          5115 => x"09",
          5116 => x"72",
          5117 => x"73",
          5118 => x"53",
          5119 => x"70",
          5120 => x"38",
          5121 => x"19",
          5122 => x"75",
          5123 => x"38",
          5124 => x"83",
          5125 => x"74",
          5126 => x"59",
          5127 => x"39",
          5128 => x"33",
          5129 => x"85",
          5130 => x"3d",
          5131 => x"3d",
          5132 => x"80",
          5133 => x"34",
          5134 => x"17",
          5135 => x"75",
          5136 => x"3f",
          5137 => x"85",
          5138 => x"82",
          5139 => x"16",
          5140 => x"3f",
          5141 => x"08",
          5142 => x"06",
          5143 => x"73",
          5144 => x"2e",
          5145 => x"80",
          5146 => x"0b",
          5147 => x"56",
          5148 => x"e9",
          5149 => x"06",
          5150 => x"57",
          5151 => x"32",
          5152 => x"05",
          5153 => x"79",
          5154 => x"54",
          5155 => x"74",
          5156 => x"09",
          5157 => x"38",
          5158 => x"fe",
          5159 => x"ea",
          5160 => x"8a",
          5161 => x"ec",
          5162 => x"85",
          5163 => x"2e",
          5164 => x"53",
          5165 => x"52",
          5166 => x"51",
          5167 => x"82",
          5168 => x"55",
          5169 => x"08",
          5170 => x"38",
          5171 => x"82",
          5172 => x"88",
          5173 => x"f1",
          5174 => x"02",
          5175 => x"cf",
          5176 => x"55",
          5177 => x"61",
          5178 => x"3f",
          5179 => x"08",
          5180 => x"80",
          5181 => x"ec",
          5182 => x"83",
          5183 => x"ec",
          5184 => x"82",
          5185 => x"08",
          5186 => x"56",
          5187 => x"86",
          5188 => x"75",
          5189 => x"fe",
          5190 => x"54",
          5191 => x"2e",
          5192 => x"14",
          5193 => x"a4",
          5194 => x"ec",
          5195 => x"06",
          5196 => x"54",
          5197 => x"38",
          5198 => x"86",
          5199 => x"82",
          5200 => x"06",
          5201 => x"56",
          5202 => x"38",
          5203 => x"80",
          5204 => x"81",
          5205 => x"52",
          5206 => x"51",
          5207 => x"82",
          5208 => x"81",
          5209 => x"81",
          5210 => x"83",
          5211 => x"8f",
          5212 => x"2e",
          5213 => x"82",
          5214 => x"06",
          5215 => x"56",
          5216 => x"38",
          5217 => x"74",
          5218 => x"a2",
          5219 => x"ec",
          5220 => x"06",
          5221 => x"2e",
          5222 => x"80",
          5223 => x"3d",
          5224 => x"83",
          5225 => x"15",
          5226 => x"53",
          5227 => x"8d",
          5228 => x"15",
          5229 => x"3f",
          5230 => x"08",
          5231 => x"70",
          5232 => x"0c",
          5233 => x"16",
          5234 => x"80",
          5235 => x"80",
          5236 => x"54",
          5237 => x"84",
          5238 => x"5c",
          5239 => x"80",
          5240 => x"7b",
          5241 => x"fc",
          5242 => x"85",
          5243 => x"ff",
          5244 => x"77",
          5245 => x"81",
          5246 => x"76",
          5247 => x"81",
          5248 => x"2e",
          5249 => x"8d",
          5250 => x"26",
          5251 => x"bf",
          5252 => x"ce",
          5253 => x"ec",
          5254 => x"ff",
          5255 => x"84",
          5256 => x"81",
          5257 => x"38",
          5258 => x"51",
          5259 => x"82",
          5260 => x"83",
          5261 => x"58",
          5262 => x"80",
          5263 => x"db",
          5264 => x"85",
          5265 => x"77",
          5266 => x"80",
          5267 => x"82",
          5268 => x"c4",
          5269 => x"11",
          5270 => x"06",
          5271 => x"8d",
          5272 => x"26",
          5273 => x"74",
          5274 => x"52",
          5275 => x"f8",
          5276 => x"85",
          5277 => x"c1",
          5278 => x"58",
          5279 => x"23",
          5280 => x"8b",
          5281 => x"73",
          5282 => x"80",
          5283 => x"8d",
          5284 => x"39",
          5285 => x"51",
          5286 => x"82",
          5287 => x"53",
          5288 => x"08",
          5289 => x"72",
          5290 => x"8d",
          5291 => x"cf",
          5292 => x"14",
          5293 => x"3f",
          5294 => x"08",
          5295 => x"06",
          5296 => x"38",
          5297 => x"51",
          5298 => x"82",
          5299 => x"55",
          5300 => x"51",
          5301 => x"82",
          5302 => x"83",
          5303 => x"5a",
          5304 => x"80",
          5305 => x"38",
          5306 => x"78",
          5307 => x"2a",
          5308 => x"78",
          5309 => x"87",
          5310 => x"22",
          5311 => x"31",
          5312 => x"87",
          5313 => x"ec",
          5314 => x"85",
          5315 => x"2e",
          5316 => x"82",
          5317 => x"80",
          5318 => x"f5",
          5319 => x"83",
          5320 => x"ff",
          5321 => x"38",
          5322 => x"9f",
          5323 => x"38",
          5324 => x"39",
          5325 => x"80",
          5326 => x"38",
          5327 => x"98",
          5328 => x"a0",
          5329 => x"1d",
          5330 => x"0c",
          5331 => x"17",
          5332 => x"76",
          5333 => x"81",
          5334 => x"80",
          5335 => x"d9",
          5336 => x"85",
          5337 => x"ff",
          5338 => x"8d",
          5339 => x"8f",
          5340 => x"8b",
          5341 => x"14",
          5342 => x"3f",
          5343 => x"08",
          5344 => x"74",
          5345 => x"a3",
          5346 => x"7a",
          5347 => x"ef",
          5348 => x"a8",
          5349 => x"15",
          5350 => x"2e",
          5351 => x"10",
          5352 => x"2a",
          5353 => x"11",
          5354 => x"83",
          5355 => x"2a",
          5356 => x"72",
          5357 => x"26",
          5358 => x"ff",
          5359 => x"0c",
          5360 => x"15",
          5361 => x"0b",
          5362 => x"76",
          5363 => x"81",
          5364 => x"38",
          5365 => x"51",
          5366 => x"82",
          5367 => x"83",
          5368 => x"53",
          5369 => x"09",
          5370 => x"f9",
          5371 => x"52",
          5372 => x"8a",
          5373 => x"ec",
          5374 => x"38",
          5375 => x"08",
          5376 => x"84",
          5377 => x"d7",
          5378 => x"85",
          5379 => x"ff",
          5380 => x"72",
          5381 => x"2e",
          5382 => x"80",
          5383 => x"14",
          5384 => x"3f",
          5385 => x"08",
          5386 => x"a4",
          5387 => x"81",
          5388 => x"84",
          5389 => x"d7",
          5390 => x"85",
          5391 => x"8a",
          5392 => x"2e",
          5393 => x"9d",
          5394 => x"14",
          5395 => x"3f",
          5396 => x"08",
          5397 => x"84",
          5398 => x"d7",
          5399 => x"85",
          5400 => x"15",
          5401 => x"34",
          5402 => x"22",
          5403 => x"72",
          5404 => x"23",
          5405 => x"23",
          5406 => x"15",
          5407 => x"75",
          5408 => x"0c",
          5409 => x"04",
          5410 => x"77",
          5411 => x"73",
          5412 => x"38",
          5413 => x"72",
          5414 => x"38",
          5415 => x"71",
          5416 => x"38",
          5417 => x"84",
          5418 => x"52",
          5419 => x"09",
          5420 => x"38",
          5421 => x"51",
          5422 => x"82",
          5423 => x"81",
          5424 => x"88",
          5425 => x"08",
          5426 => x"39",
          5427 => x"73",
          5428 => x"74",
          5429 => x"0c",
          5430 => x"04",
          5431 => x"02",
          5432 => x"7a",
          5433 => x"fc",
          5434 => x"f4",
          5435 => x"54",
          5436 => x"85",
          5437 => x"bc",
          5438 => x"ec",
          5439 => x"82",
          5440 => x"70",
          5441 => x"73",
          5442 => x"38",
          5443 => x"78",
          5444 => x"2e",
          5445 => x"74",
          5446 => x"0c",
          5447 => x"80",
          5448 => x"80",
          5449 => x"70",
          5450 => x"51",
          5451 => x"82",
          5452 => x"54",
          5453 => x"ec",
          5454 => x"0d",
          5455 => x"0d",
          5456 => x"05",
          5457 => x"33",
          5458 => x"54",
          5459 => x"84",
          5460 => x"bf",
          5461 => x"98",
          5462 => x"53",
          5463 => x"05",
          5464 => x"f3",
          5465 => x"ec",
          5466 => x"85",
          5467 => x"a6",
          5468 => x"68",
          5469 => x"70",
          5470 => x"a7",
          5471 => x"ec",
          5472 => x"85",
          5473 => x"38",
          5474 => x"05",
          5475 => x"2b",
          5476 => x"80",
          5477 => x"86",
          5478 => x"06",
          5479 => x"2e",
          5480 => x"74",
          5481 => x"38",
          5482 => x"09",
          5483 => x"38",
          5484 => x"d9",
          5485 => x"ec",
          5486 => x"39",
          5487 => x"33",
          5488 => x"73",
          5489 => x"77",
          5490 => x"81",
          5491 => x"73",
          5492 => x"38",
          5493 => x"be",
          5494 => x"07",
          5495 => x"b6",
          5496 => x"2a",
          5497 => x"51",
          5498 => x"2e",
          5499 => x"62",
          5500 => x"e8",
          5501 => x"85",
          5502 => x"82",
          5503 => x"52",
          5504 => x"51",
          5505 => x"62",
          5506 => x"8b",
          5507 => x"53",
          5508 => x"51",
          5509 => x"80",
          5510 => x"05",
          5511 => x"3f",
          5512 => x"0b",
          5513 => x"75",
          5514 => x"f1",
          5515 => x"11",
          5516 => x"80",
          5517 => x"97",
          5518 => x"51",
          5519 => x"82",
          5520 => x"55",
          5521 => x"08",
          5522 => x"b7",
          5523 => x"c6",
          5524 => x"05",
          5525 => x"2a",
          5526 => x"51",
          5527 => x"80",
          5528 => x"84",
          5529 => x"39",
          5530 => x"70",
          5531 => x"54",
          5532 => x"a9",
          5533 => x"06",
          5534 => x"2e",
          5535 => x"55",
          5536 => x"73",
          5537 => x"d5",
          5538 => x"85",
          5539 => x"ff",
          5540 => x"0c",
          5541 => x"85",
          5542 => x"fa",
          5543 => x"2a",
          5544 => x"51",
          5545 => x"2e",
          5546 => x"80",
          5547 => x"7a",
          5548 => x"a0",
          5549 => x"a4",
          5550 => x"53",
          5551 => x"e6",
          5552 => x"85",
          5553 => x"85",
          5554 => x"1b",
          5555 => x"05",
          5556 => x"a5",
          5557 => x"ec",
          5558 => x"ec",
          5559 => x"0c",
          5560 => x"56",
          5561 => x"84",
          5562 => x"90",
          5563 => x"0b",
          5564 => x"80",
          5565 => x"0c",
          5566 => x"1a",
          5567 => x"2a",
          5568 => x"51",
          5569 => x"2e",
          5570 => x"82",
          5571 => x"80",
          5572 => x"38",
          5573 => x"08",
          5574 => x"8a",
          5575 => x"89",
          5576 => x"59",
          5577 => x"76",
          5578 => x"d6",
          5579 => x"85",
          5580 => x"82",
          5581 => x"81",
          5582 => x"82",
          5583 => x"ec",
          5584 => x"09",
          5585 => x"38",
          5586 => x"78",
          5587 => x"09",
          5588 => x"76",
          5589 => x"51",
          5590 => x"27",
          5591 => x"70",
          5592 => x"5a",
          5593 => x"76",
          5594 => x"74",
          5595 => x"83",
          5596 => x"73",
          5597 => x"38",
          5598 => x"51",
          5599 => x"82",
          5600 => x"85",
          5601 => x"8e",
          5602 => x"2a",
          5603 => x"08",
          5604 => x"0c",
          5605 => x"79",
          5606 => x"73",
          5607 => x"0c",
          5608 => x"04",
          5609 => x"60",
          5610 => x"40",
          5611 => x"80",
          5612 => x"3d",
          5613 => x"78",
          5614 => x"3f",
          5615 => x"08",
          5616 => x"ec",
          5617 => x"91",
          5618 => x"74",
          5619 => x"38",
          5620 => x"c4",
          5621 => x"33",
          5622 => x"87",
          5623 => x"2e",
          5624 => x"95",
          5625 => x"91",
          5626 => x"56",
          5627 => x"81",
          5628 => x"34",
          5629 => x"a0",
          5630 => x"08",
          5631 => x"31",
          5632 => x"27",
          5633 => x"5c",
          5634 => x"82",
          5635 => x"19",
          5636 => x"ff",
          5637 => x"74",
          5638 => x"7e",
          5639 => x"ff",
          5640 => x"2a",
          5641 => x"79",
          5642 => x"87",
          5643 => x"08",
          5644 => x"98",
          5645 => x"78",
          5646 => x"3f",
          5647 => x"08",
          5648 => x"27",
          5649 => x"74",
          5650 => x"a3",
          5651 => x"1a",
          5652 => x"08",
          5653 => x"d4",
          5654 => x"85",
          5655 => x"2e",
          5656 => x"82",
          5657 => x"1a",
          5658 => x"59",
          5659 => x"2e",
          5660 => x"77",
          5661 => x"11",
          5662 => x"55",
          5663 => x"85",
          5664 => x"31",
          5665 => x"76",
          5666 => x"81",
          5667 => x"c9",
          5668 => x"85",
          5669 => x"d7",
          5670 => x"11",
          5671 => x"74",
          5672 => x"38",
          5673 => x"77",
          5674 => x"78",
          5675 => x"84",
          5676 => x"16",
          5677 => x"08",
          5678 => x"2b",
          5679 => x"cf",
          5680 => x"89",
          5681 => x"39",
          5682 => x"0c",
          5683 => x"83",
          5684 => x"80",
          5685 => x"55",
          5686 => x"83",
          5687 => x"9c",
          5688 => x"7e",
          5689 => x"3f",
          5690 => x"08",
          5691 => x"75",
          5692 => x"08",
          5693 => x"1f",
          5694 => x"7c",
          5695 => x"3f",
          5696 => x"7e",
          5697 => x"0c",
          5698 => x"1b",
          5699 => x"1c",
          5700 => x"fd",
          5701 => x"56",
          5702 => x"ec",
          5703 => x"0d",
          5704 => x"0d",
          5705 => x"64",
          5706 => x"58",
          5707 => x"90",
          5708 => x"52",
          5709 => x"d0",
          5710 => x"ec",
          5711 => x"85",
          5712 => x"38",
          5713 => x"55",
          5714 => x"86",
          5715 => x"83",
          5716 => x"18",
          5717 => x"2a",
          5718 => x"51",
          5719 => x"56",
          5720 => x"83",
          5721 => x"39",
          5722 => x"19",
          5723 => x"83",
          5724 => x"0b",
          5725 => x"81",
          5726 => x"39",
          5727 => x"7c",
          5728 => x"74",
          5729 => x"38",
          5730 => x"7b",
          5731 => x"ec",
          5732 => x"08",
          5733 => x"06",
          5734 => x"81",
          5735 => x"8a",
          5736 => x"05",
          5737 => x"06",
          5738 => x"bf",
          5739 => x"38",
          5740 => x"55",
          5741 => x"7a",
          5742 => x"98",
          5743 => x"77",
          5744 => x"3f",
          5745 => x"08",
          5746 => x"ec",
          5747 => x"82",
          5748 => x"81",
          5749 => x"38",
          5750 => x"ff",
          5751 => x"98",
          5752 => x"18",
          5753 => x"74",
          5754 => x"7e",
          5755 => x"08",
          5756 => x"2e",
          5757 => x"8d",
          5758 => x"ce",
          5759 => x"85",
          5760 => x"ee",
          5761 => x"08",
          5762 => x"d0",
          5763 => x"85",
          5764 => x"2e",
          5765 => x"82",
          5766 => x"1b",
          5767 => x"5a",
          5768 => x"2e",
          5769 => x"78",
          5770 => x"11",
          5771 => x"55",
          5772 => x"85",
          5773 => x"31",
          5774 => x"76",
          5775 => x"81",
          5776 => x"c8",
          5777 => x"85",
          5778 => x"a6",
          5779 => x"11",
          5780 => x"56",
          5781 => x"27",
          5782 => x"80",
          5783 => x"08",
          5784 => x"2b",
          5785 => x"b4",
          5786 => x"85",
          5787 => x"80",
          5788 => x"34",
          5789 => x"56",
          5790 => x"8c",
          5791 => x"19",
          5792 => x"38",
          5793 => x"86",
          5794 => x"ec",
          5795 => x"38",
          5796 => x"12",
          5797 => x"9c",
          5798 => x"18",
          5799 => x"06",
          5800 => x"31",
          5801 => x"76",
          5802 => x"7b",
          5803 => x"08",
          5804 => x"cd",
          5805 => x"85",
          5806 => x"b6",
          5807 => x"7c",
          5808 => x"08",
          5809 => x"1f",
          5810 => x"cb",
          5811 => x"55",
          5812 => x"16",
          5813 => x"31",
          5814 => x"7f",
          5815 => x"94",
          5816 => x"70",
          5817 => x"8c",
          5818 => x"58",
          5819 => x"76",
          5820 => x"75",
          5821 => x"19",
          5822 => x"39",
          5823 => x"80",
          5824 => x"74",
          5825 => x"80",
          5826 => x"85",
          5827 => x"3d",
          5828 => x"3d",
          5829 => x"3d",
          5830 => x"70",
          5831 => x"e8",
          5832 => x"ec",
          5833 => x"85",
          5834 => x"fb",
          5835 => x"33",
          5836 => x"70",
          5837 => x"55",
          5838 => x"2e",
          5839 => x"a0",
          5840 => x"78",
          5841 => x"3f",
          5842 => x"08",
          5843 => x"ec",
          5844 => x"38",
          5845 => x"8b",
          5846 => x"07",
          5847 => x"8b",
          5848 => x"16",
          5849 => x"52",
          5850 => x"dd",
          5851 => x"16",
          5852 => x"15",
          5853 => x"3f",
          5854 => x"0a",
          5855 => x"51",
          5856 => x"76",
          5857 => x"51",
          5858 => x"78",
          5859 => x"83",
          5860 => x"51",
          5861 => x"82",
          5862 => x"90",
          5863 => x"bf",
          5864 => x"73",
          5865 => x"76",
          5866 => x"0c",
          5867 => x"04",
          5868 => x"76",
          5869 => x"fe",
          5870 => x"85",
          5871 => x"82",
          5872 => x"9c",
          5873 => x"fc",
          5874 => x"51",
          5875 => x"82",
          5876 => x"53",
          5877 => x"08",
          5878 => x"85",
          5879 => x"0c",
          5880 => x"ec",
          5881 => x"0d",
          5882 => x"0d",
          5883 => x"e6",
          5884 => x"52",
          5885 => x"85",
          5886 => x"8b",
          5887 => x"ec",
          5888 => x"a4",
          5889 => x"71",
          5890 => x"0c",
          5891 => x"04",
          5892 => x"80",
          5893 => x"d0",
          5894 => x"3d",
          5895 => x"3f",
          5896 => x"08",
          5897 => x"ec",
          5898 => x"38",
          5899 => x"52",
          5900 => x"05",
          5901 => x"3f",
          5902 => x"08",
          5903 => x"ec",
          5904 => x"02",
          5905 => x"33",
          5906 => x"55",
          5907 => x"25",
          5908 => x"7a",
          5909 => x"54",
          5910 => x"a2",
          5911 => x"84",
          5912 => x"06",
          5913 => x"73",
          5914 => x"38",
          5915 => x"70",
          5916 => x"87",
          5917 => x"ec",
          5918 => x"0c",
          5919 => x"85",
          5920 => x"2e",
          5921 => x"83",
          5922 => x"74",
          5923 => x"0c",
          5924 => x"04",
          5925 => x"6f",
          5926 => x"80",
          5927 => x"53",
          5928 => x"b8",
          5929 => x"3d",
          5930 => x"3f",
          5931 => x"08",
          5932 => x"ec",
          5933 => x"38",
          5934 => x"7c",
          5935 => x"47",
          5936 => x"54",
          5937 => x"81",
          5938 => x"52",
          5939 => x"52",
          5940 => x"3f",
          5941 => x"08",
          5942 => x"ec",
          5943 => x"38",
          5944 => x"51",
          5945 => x"82",
          5946 => x"57",
          5947 => x"08",
          5948 => x"69",
          5949 => x"da",
          5950 => x"85",
          5951 => x"76",
          5952 => x"d5",
          5953 => x"85",
          5954 => x"82",
          5955 => x"82",
          5956 => x"52",
          5957 => x"ca",
          5958 => x"ec",
          5959 => x"85",
          5960 => x"38",
          5961 => x"51",
          5962 => x"73",
          5963 => x"08",
          5964 => x"76",
          5965 => x"d6",
          5966 => x"85",
          5967 => x"82",
          5968 => x"80",
          5969 => x"76",
          5970 => x"81",
          5971 => x"82",
          5972 => x"39",
          5973 => x"38",
          5974 => x"bc",
          5975 => x"51",
          5976 => x"76",
          5977 => x"11",
          5978 => x"51",
          5979 => x"73",
          5980 => x"38",
          5981 => x"55",
          5982 => x"16",
          5983 => x"56",
          5984 => x"38",
          5985 => x"73",
          5986 => x"8f",
          5987 => x"2e",
          5988 => x"16",
          5989 => x"ff",
          5990 => x"ff",
          5991 => x"58",
          5992 => x"74",
          5993 => x"75",
          5994 => x"18",
          5995 => x"58",
          5996 => x"fe",
          5997 => x"7b",
          5998 => x"06",
          5999 => x"18",
          6000 => x"58",
          6001 => x"80",
          6002 => x"a4",
          6003 => x"2b",
          6004 => x"11",
          6005 => x"52",
          6006 => x"56",
          6007 => x"8d",
          6008 => x"70",
          6009 => x"51",
          6010 => x"f5",
          6011 => x"54",
          6012 => x"a7",
          6013 => x"74",
          6014 => x"38",
          6015 => x"73",
          6016 => x"81",
          6017 => x"81",
          6018 => x"39",
          6019 => x"81",
          6020 => x"74",
          6021 => x"81",
          6022 => x"91",
          6023 => x"6e",
          6024 => x"59",
          6025 => x"7a",
          6026 => x"5c",
          6027 => x"26",
          6028 => x"7a",
          6029 => x"85",
          6030 => x"3d",
          6031 => x"3d",
          6032 => x"8d",
          6033 => x"54",
          6034 => x"55",
          6035 => x"82",
          6036 => x"53",
          6037 => x"08",
          6038 => x"91",
          6039 => x"72",
          6040 => x"8c",
          6041 => x"73",
          6042 => x"38",
          6043 => x"70",
          6044 => x"81",
          6045 => x"57",
          6046 => x"73",
          6047 => x"08",
          6048 => x"94",
          6049 => x"75",
          6050 => x"99",
          6051 => x"11",
          6052 => x"2b",
          6053 => x"73",
          6054 => x"38",
          6055 => x"16",
          6056 => x"e7",
          6057 => x"ec",
          6058 => x"78",
          6059 => x"55",
          6060 => x"d7",
          6061 => x"ec",
          6062 => x"98",
          6063 => x"81",
          6064 => x"06",
          6065 => x"0c",
          6066 => x"98",
          6067 => x"58",
          6068 => x"39",
          6069 => x"54",
          6070 => x"73",
          6071 => x"cd",
          6072 => x"85",
          6073 => x"82",
          6074 => x"81",
          6075 => x"38",
          6076 => x"08",
          6077 => x"9b",
          6078 => x"ec",
          6079 => x"0c",
          6080 => x"0c",
          6081 => x"81",
          6082 => x"76",
          6083 => x"38",
          6084 => x"94",
          6085 => x"94",
          6086 => x"16",
          6087 => x"2a",
          6088 => x"51",
          6089 => x"72",
          6090 => x"38",
          6091 => x"51",
          6092 => x"82",
          6093 => x"54",
          6094 => x"08",
          6095 => x"85",
          6096 => x"a7",
          6097 => x"74",
          6098 => x"3f",
          6099 => x"08",
          6100 => x"2e",
          6101 => x"74",
          6102 => x"79",
          6103 => x"14",
          6104 => x"38",
          6105 => x"0c",
          6106 => x"94",
          6107 => x"94",
          6108 => x"83",
          6109 => x"72",
          6110 => x"38",
          6111 => x"51",
          6112 => x"82",
          6113 => x"94",
          6114 => x"91",
          6115 => x"53",
          6116 => x"81",
          6117 => x"34",
          6118 => x"39",
          6119 => x"82",
          6120 => x"05",
          6121 => x"08",
          6122 => x"08",
          6123 => x"38",
          6124 => x"0c",
          6125 => x"80",
          6126 => x"72",
          6127 => x"73",
          6128 => x"53",
          6129 => x"8c",
          6130 => x"16",
          6131 => x"38",
          6132 => x"0c",
          6133 => x"82",
          6134 => x"8b",
          6135 => x"f9",
          6136 => x"56",
          6137 => x"80",
          6138 => x"38",
          6139 => x"3d",
          6140 => x"8a",
          6141 => x"51",
          6142 => x"82",
          6143 => x"55",
          6144 => x"08",
          6145 => x"77",
          6146 => x"52",
          6147 => x"93",
          6148 => x"ec",
          6149 => x"85",
          6150 => x"c3",
          6151 => x"33",
          6152 => x"55",
          6153 => x"24",
          6154 => x"16",
          6155 => x"2a",
          6156 => x"51",
          6157 => x"80",
          6158 => x"9c",
          6159 => x"77",
          6160 => x"3f",
          6161 => x"08",
          6162 => x"77",
          6163 => x"22",
          6164 => x"74",
          6165 => x"ce",
          6166 => x"85",
          6167 => x"74",
          6168 => x"81",
          6169 => x"85",
          6170 => x"74",
          6171 => x"38",
          6172 => x"74",
          6173 => x"85",
          6174 => x"3d",
          6175 => x"3d",
          6176 => x"3d",
          6177 => x"70",
          6178 => x"fc",
          6179 => x"ec",
          6180 => x"82",
          6181 => x"73",
          6182 => x"0d",
          6183 => x"0d",
          6184 => x"3d",
          6185 => x"71",
          6186 => x"e7",
          6187 => x"85",
          6188 => x"82",
          6189 => x"80",
          6190 => x"93",
          6191 => x"ec",
          6192 => x"51",
          6193 => x"82",
          6194 => x"53",
          6195 => x"82",
          6196 => x"52",
          6197 => x"8a",
          6198 => x"ec",
          6199 => x"85",
          6200 => x"2e",
          6201 => x"85",
          6202 => x"87",
          6203 => x"ec",
          6204 => x"74",
          6205 => x"d5",
          6206 => x"52",
          6207 => x"e7",
          6208 => x"ec",
          6209 => x"70",
          6210 => x"70",
          6211 => x"2c",
          6212 => x"ec",
          6213 => x"51",
          6214 => x"82",
          6215 => x"87",
          6216 => x"ee",
          6217 => x"57",
          6218 => x"3d",
          6219 => x"3d",
          6220 => x"a3",
          6221 => x"ec",
          6222 => x"85",
          6223 => x"38",
          6224 => x"51",
          6225 => x"82",
          6226 => x"55",
          6227 => x"08",
          6228 => x"80",
          6229 => x"70",
          6230 => x"58",
          6231 => x"85",
          6232 => x"8d",
          6233 => x"2e",
          6234 => x"52",
          6235 => x"9a",
          6236 => x"85",
          6237 => x"3d",
          6238 => x"3d",
          6239 => x"55",
          6240 => x"92",
          6241 => x"52",
          6242 => x"de",
          6243 => x"85",
          6244 => x"82",
          6245 => x"82",
          6246 => x"74",
          6247 => x"98",
          6248 => x"11",
          6249 => x"59",
          6250 => x"75",
          6251 => x"38",
          6252 => x"81",
          6253 => x"5b",
          6254 => x"82",
          6255 => x"39",
          6256 => x"08",
          6257 => x"59",
          6258 => x"09",
          6259 => x"c1",
          6260 => x"5f",
          6261 => x"92",
          6262 => x"51",
          6263 => x"82",
          6264 => x"ff",
          6265 => x"82",
          6266 => x"81",
          6267 => x"82",
          6268 => x"09",
          6269 => x"82",
          6270 => x"07",
          6271 => x"05",
          6272 => x"53",
          6273 => x"98",
          6274 => x"26",
          6275 => x"fd",
          6276 => x"08",
          6277 => x"08",
          6278 => x"98",
          6279 => x"81",
          6280 => x"58",
          6281 => x"3f",
          6282 => x"08",
          6283 => x"ec",
          6284 => x"38",
          6285 => x"77",
          6286 => x"5d",
          6287 => x"74",
          6288 => x"81",
          6289 => x"b4",
          6290 => x"bb",
          6291 => x"85",
          6292 => x"ff",
          6293 => x"09",
          6294 => x"80",
          6295 => x"19",
          6296 => x"54",
          6297 => x"14",
          6298 => x"8d",
          6299 => x"ec",
          6300 => x"06",
          6301 => x"05",
          6302 => x"1b",
          6303 => x"5b",
          6304 => x"83",
          6305 => x"58",
          6306 => x"8e",
          6307 => x"0c",
          6308 => x"12",
          6309 => x"33",
          6310 => x"54",
          6311 => x"34",
          6312 => x"ec",
          6313 => x"0d",
          6314 => x"0d",
          6315 => x"fc",
          6316 => x"52",
          6317 => x"3f",
          6318 => x"08",
          6319 => x"ec",
          6320 => x"38",
          6321 => x"56",
          6322 => x"38",
          6323 => x"70",
          6324 => x"81",
          6325 => x"55",
          6326 => x"80",
          6327 => x"38",
          6328 => x"54",
          6329 => x"08",
          6330 => x"38",
          6331 => x"82",
          6332 => x"53",
          6333 => x"52",
          6334 => x"d9",
          6335 => x"ec",
          6336 => x"19",
          6337 => x"c9",
          6338 => x"08",
          6339 => x"ff",
          6340 => x"82",
          6341 => x"ff",
          6342 => x"06",
          6343 => x"56",
          6344 => x"08",
          6345 => x"81",
          6346 => x"82",
          6347 => x"75",
          6348 => x"54",
          6349 => x"08",
          6350 => x"27",
          6351 => x"17",
          6352 => x"85",
          6353 => x"76",
          6354 => x"3f",
          6355 => x"08",
          6356 => x"08",
          6357 => x"90",
          6358 => x"c0",
          6359 => x"90",
          6360 => x"80",
          6361 => x"75",
          6362 => x"75",
          6363 => x"85",
          6364 => x"3d",
          6365 => x"3d",
          6366 => x"a0",
          6367 => x"05",
          6368 => x"51",
          6369 => x"82",
          6370 => x"55",
          6371 => x"08",
          6372 => x"78",
          6373 => x"08",
          6374 => x"70",
          6375 => x"83",
          6376 => x"ec",
          6377 => x"85",
          6378 => x"dd",
          6379 => x"fb",
          6380 => x"85",
          6381 => x"06",
          6382 => x"86",
          6383 => x"c9",
          6384 => x"2b",
          6385 => x"24",
          6386 => x"02",
          6387 => x"33",
          6388 => x"58",
          6389 => x"76",
          6390 => x"6b",
          6391 => x"cc",
          6392 => x"85",
          6393 => x"84",
          6394 => x"06",
          6395 => x"73",
          6396 => x"d4",
          6397 => x"82",
          6398 => x"94",
          6399 => x"81",
          6400 => x"5a",
          6401 => x"08",
          6402 => x"8a",
          6403 => x"54",
          6404 => x"82",
          6405 => x"55",
          6406 => x"08",
          6407 => x"82",
          6408 => x"52",
          6409 => x"ba",
          6410 => x"ec",
          6411 => x"85",
          6412 => x"38",
          6413 => x"d1",
          6414 => x"ec",
          6415 => x"88",
          6416 => x"ec",
          6417 => x"38",
          6418 => x"97",
          6419 => x"ec",
          6420 => x"ec",
          6421 => x"05",
          6422 => x"ec",
          6423 => x"25",
          6424 => x"75",
          6425 => x"38",
          6426 => x"8f",
          6427 => x"75",
          6428 => x"c0",
          6429 => x"85",
          6430 => x"74",
          6431 => x"51",
          6432 => x"3f",
          6433 => x"08",
          6434 => x"85",
          6435 => x"3d",
          6436 => x"3d",
          6437 => x"99",
          6438 => x"52",
          6439 => x"d8",
          6440 => x"85",
          6441 => x"82",
          6442 => x"82",
          6443 => x"5e",
          6444 => x"3d",
          6445 => x"ce",
          6446 => x"85",
          6447 => x"82",
          6448 => x"86",
          6449 => x"82",
          6450 => x"85",
          6451 => x"2e",
          6452 => x"82",
          6453 => x"80",
          6454 => x"70",
          6455 => x"06",
          6456 => x"54",
          6457 => x"38",
          6458 => x"52",
          6459 => x"52",
          6460 => x"3f",
          6461 => x"08",
          6462 => x"82",
          6463 => x"83",
          6464 => x"82",
          6465 => x"81",
          6466 => x"06",
          6467 => x"54",
          6468 => x"08",
          6469 => x"81",
          6470 => x"81",
          6471 => x"39",
          6472 => x"38",
          6473 => x"08",
          6474 => x"c3",
          6475 => x"85",
          6476 => x"82",
          6477 => x"81",
          6478 => x"53",
          6479 => x"19",
          6480 => x"d0",
          6481 => x"ae",
          6482 => x"34",
          6483 => x"0b",
          6484 => x"82",
          6485 => x"52",
          6486 => x"51",
          6487 => x"3f",
          6488 => x"b4",
          6489 => x"c9",
          6490 => x"53",
          6491 => x"53",
          6492 => x"51",
          6493 => x"3f",
          6494 => x"0b",
          6495 => x"34",
          6496 => x"80",
          6497 => x"51",
          6498 => x"78",
          6499 => x"83",
          6500 => x"51",
          6501 => x"82",
          6502 => x"54",
          6503 => x"08",
          6504 => x"88",
          6505 => x"64",
          6506 => x"ff",
          6507 => x"75",
          6508 => x"78",
          6509 => x"3f",
          6510 => x"0b",
          6511 => x"78",
          6512 => x"83",
          6513 => x"51",
          6514 => x"3f",
          6515 => x"08",
          6516 => x"80",
          6517 => x"76",
          6518 => x"f9",
          6519 => x"85",
          6520 => x"3d",
          6521 => x"3d",
          6522 => x"84",
          6523 => x"d4",
          6524 => x"a8",
          6525 => x"05",
          6526 => x"51",
          6527 => x"82",
          6528 => x"55",
          6529 => x"08",
          6530 => x"78",
          6531 => x"08",
          6532 => x"70",
          6533 => x"8b",
          6534 => x"ec",
          6535 => x"85",
          6536 => x"b9",
          6537 => x"9b",
          6538 => x"a0",
          6539 => x"55",
          6540 => x"38",
          6541 => x"3d",
          6542 => x"3d",
          6543 => x"51",
          6544 => x"3f",
          6545 => x"52",
          6546 => x"52",
          6547 => x"a1",
          6548 => x"08",
          6549 => x"cb",
          6550 => x"85",
          6551 => x"82",
          6552 => x"95",
          6553 => x"2e",
          6554 => x"88",
          6555 => x"3d",
          6556 => x"38",
          6557 => x"e5",
          6558 => x"ec",
          6559 => x"09",
          6560 => x"b8",
          6561 => x"c9",
          6562 => x"85",
          6563 => x"82",
          6564 => x"81",
          6565 => x"56",
          6566 => x"3d",
          6567 => x"52",
          6568 => x"ff",
          6569 => x"02",
          6570 => x"8b",
          6571 => x"16",
          6572 => x"2a",
          6573 => x"51",
          6574 => x"89",
          6575 => x"07",
          6576 => x"17",
          6577 => x"81",
          6578 => x"34",
          6579 => x"70",
          6580 => x"81",
          6581 => x"55",
          6582 => x"80",
          6583 => x"64",
          6584 => x"38",
          6585 => x"51",
          6586 => x"82",
          6587 => x"52",
          6588 => x"b6",
          6589 => x"55",
          6590 => x"08",
          6591 => x"dd",
          6592 => x"ec",
          6593 => x"51",
          6594 => x"3f",
          6595 => x"08",
          6596 => x"11",
          6597 => x"82",
          6598 => x"80",
          6599 => x"16",
          6600 => x"ae",
          6601 => x"06",
          6602 => x"53",
          6603 => x"51",
          6604 => x"78",
          6605 => x"83",
          6606 => x"39",
          6607 => x"08",
          6608 => x"51",
          6609 => x"82",
          6610 => x"55",
          6611 => x"08",
          6612 => x"51",
          6613 => x"3f",
          6614 => x"08",
          6615 => x"85",
          6616 => x"3d",
          6617 => x"3d",
          6618 => x"db",
          6619 => x"84",
          6620 => x"05",
          6621 => x"82",
          6622 => x"d0",
          6623 => x"3d",
          6624 => x"3f",
          6625 => x"08",
          6626 => x"ec",
          6627 => x"38",
          6628 => x"52",
          6629 => x"05",
          6630 => x"3f",
          6631 => x"08",
          6632 => x"ec",
          6633 => x"02",
          6634 => x"33",
          6635 => x"54",
          6636 => x"aa",
          6637 => x"06",
          6638 => x"8b",
          6639 => x"06",
          6640 => x"07",
          6641 => x"56",
          6642 => x"34",
          6643 => x"0b",
          6644 => x"78",
          6645 => x"ed",
          6646 => x"ec",
          6647 => x"82",
          6648 => x"95",
          6649 => x"ef",
          6650 => x"56",
          6651 => x"3d",
          6652 => x"94",
          6653 => x"df",
          6654 => x"ec",
          6655 => x"85",
          6656 => x"cb",
          6657 => x"63",
          6658 => x"d4",
          6659 => x"93",
          6660 => x"ec",
          6661 => x"85",
          6662 => x"38",
          6663 => x"05",
          6664 => x"06",
          6665 => x"73",
          6666 => x"16",
          6667 => x"22",
          6668 => x"07",
          6669 => x"1f",
          6670 => x"86",
          6671 => x"81",
          6672 => x"34",
          6673 => x"b2",
          6674 => x"85",
          6675 => x"74",
          6676 => x"0c",
          6677 => x"04",
          6678 => x"69",
          6679 => x"80",
          6680 => x"d0",
          6681 => x"3d",
          6682 => x"3f",
          6683 => x"08",
          6684 => x"08",
          6685 => x"70",
          6686 => x"08",
          6687 => x"51",
          6688 => x"80",
          6689 => x"38",
          6690 => x"06",
          6691 => x"80",
          6692 => x"38",
          6693 => x"5f",
          6694 => x"3d",
          6695 => x"ff",
          6696 => x"82",
          6697 => x"57",
          6698 => x"08",
          6699 => x"74",
          6700 => x"c3",
          6701 => x"85",
          6702 => x"82",
          6703 => x"bf",
          6704 => x"ec",
          6705 => x"ec",
          6706 => x"59",
          6707 => x"81",
          6708 => x"56",
          6709 => x"33",
          6710 => x"16",
          6711 => x"27",
          6712 => x"56",
          6713 => x"80",
          6714 => x"80",
          6715 => x"ff",
          6716 => x"70",
          6717 => x"56",
          6718 => x"e8",
          6719 => x"76",
          6720 => x"81",
          6721 => x"80",
          6722 => x"57",
          6723 => x"05",
          6724 => x"80",
          6725 => x"7a",
          6726 => x"c1",
          6727 => x"2e",
          6728 => x"a0",
          6729 => x"51",
          6730 => x"3f",
          6731 => x"08",
          6732 => x"ec",
          6733 => x"7b",
          6734 => x"55",
          6735 => x"73",
          6736 => x"38",
          6737 => x"73",
          6738 => x"38",
          6739 => x"15",
          6740 => x"ff",
          6741 => x"82",
          6742 => x"7b",
          6743 => x"85",
          6744 => x"3d",
          6745 => x"3d",
          6746 => x"9c",
          6747 => x"05",
          6748 => x"51",
          6749 => x"82",
          6750 => x"82",
          6751 => x"56",
          6752 => x"ec",
          6753 => x"38",
          6754 => x"52",
          6755 => x"52",
          6756 => x"80",
          6757 => x"70",
          6758 => x"ff",
          6759 => x"55",
          6760 => x"27",
          6761 => x"78",
          6762 => x"ff",
          6763 => x"05",
          6764 => x"55",
          6765 => x"3f",
          6766 => x"08",
          6767 => x"38",
          6768 => x"70",
          6769 => x"ff",
          6770 => x"82",
          6771 => x"80",
          6772 => x"74",
          6773 => x"07",
          6774 => x"4e",
          6775 => x"82",
          6776 => x"55",
          6777 => x"70",
          6778 => x"06",
          6779 => x"99",
          6780 => x"e0",
          6781 => x"ff",
          6782 => x"54",
          6783 => x"27",
          6784 => x"fe",
          6785 => x"55",
          6786 => x"a3",
          6787 => x"82",
          6788 => x"ff",
          6789 => x"82",
          6790 => x"93",
          6791 => x"75",
          6792 => x"76",
          6793 => x"38",
          6794 => x"77",
          6795 => x"86",
          6796 => x"39",
          6797 => x"27",
          6798 => x"88",
          6799 => x"78",
          6800 => x"5a",
          6801 => x"57",
          6802 => x"81",
          6803 => x"81",
          6804 => x"33",
          6805 => x"06",
          6806 => x"57",
          6807 => x"fe",
          6808 => x"3d",
          6809 => x"55",
          6810 => x"2e",
          6811 => x"76",
          6812 => x"38",
          6813 => x"55",
          6814 => x"33",
          6815 => x"a0",
          6816 => x"06",
          6817 => x"17",
          6818 => x"38",
          6819 => x"43",
          6820 => x"3d",
          6821 => x"ff",
          6822 => x"82",
          6823 => x"54",
          6824 => x"08",
          6825 => x"81",
          6826 => x"ff",
          6827 => x"82",
          6828 => x"54",
          6829 => x"08",
          6830 => x"80",
          6831 => x"54",
          6832 => x"80",
          6833 => x"85",
          6834 => x"2e",
          6835 => x"80",
          6836 => x"54",
          6837 => x"80",
          6838 => x"52",
          6839 => x"bc",
          6840 => x"85",
          6841 => x"82",
          6842 => x"b1",
          6843 => x"82",
          6844 => x"52",
          6845 => x"ab",
          6846 => x"54",
          6847 => x"15",
          6848 => x"78",
          6849 => x"ff",
          6850 => x"79",
          6851 => x"83",
          6852 => x"51",
          6853 => x"3f",
          6854 => x"08",
          6855 => x"74",
          6856 => x"0c",
          6857 => x"04",
          6858 => x"60",
          6859 => x"05",
          6860 => x"33",
          6861 => x"05",
          6862 => x"40",
          6863 => x"c8",
          6864 => x"ec",
          6865 => x"85",
          6866 => x"bf",
          6867 => x"33",
          6868 => x"b7",
          6869 => x"2e",
          6870 => x"1a",
          6871 => x"90",
          6872 => x"33",
          6873 => x"70",
          6874 => x"55",
          6875 => x"38",
          6876 => x"99",
          6877 => x"82",
          6878 => x"58",
          6879 => x"7e",
          6880 => x"70",
          6881 => x"55",
          6882 => x"56",
          6883 => x"fb",
          6884 => x"7d",
          6885 => x"81",
          6886 => x"07",
          6887 => x"85",
          6888 => x"8c",
          6889 => x"40",
          6890 => x"55",
          6891 => x"88",
          6892 => x"08",
          6893 => x"38",
          6894 => x"77",
          6895 => x"56",
          6896 => x"51",
          6897 => x"3f",
          6898 => x"55",
          6899 => x"08",
          6900 => x"38",
          6901 => x"85",
          6902 => x"2e",
          6903 => x"82",
          6904 => x"ff",
          6905 => x"38",
          6906 => x"08",
          6907 => x"16",
          6908 => x"2e",
          6909 => x"87",
          6910 => x"74",
          6911 => x"74",
          6912 => x"81",
          6913 => x"38",
          6914 => x"ff",
          6915 => x"2e",
          6916 => x"7b",
          6917 => x"80",
          6918 => x"81",
          6919 => x"81",
          6920 => x"06",
          6921 => x"56",
          6922 => x"52",
          6923 => x"ae",
          6924 => x"85",
          6925 => x"82",
          6926 => x"80",
          6927 => x"81",
          6928 => x"56",
          6929 => x"d3",
          6930 => x"ff",
          6931 => x"7c",
          6932 => x"55",
          6933 => x"b3",
          6934 => x"1b",
          6935 => x"1b",
          6936 => x"33",
          6937 => x"54",
          6938 => x"34",
          6939 => x"fe",
          6940 => x"08",
          6941 => x"74",
          6942 => x"75",
          6943 => x"16",
          6944 => x"33",
          6945 => x"73",
          6946 => x"77",
          6947 => x"85",
          6948 => x"3d",
          6949 => x"3d",
          6950 => x"02",
          6951 => x"eb",
          6952 => x"3d",
          6953 => x"59",
          6954 => x"8b",
          6955 => x"82",
          6956 => x"24",
          6957 => x"82",
          6958 => x"82",
          6959 => x"90",
          6960 => x"55",
          6961 => x"84",
          6962 => x"34",
          6963 => x"08",
          6964 => x"5f",
          6965 => x"51",
          6966 => x"3f",
          6967 => x"08",
          6968 => x"70",
          6969 => x"57",
          6970 => x"8b",
          6971 => x"82",
          6972 => x"06",
          6973 => x"56",
          6974 => x"38",
          6975 => x"05",
          6976 => x"7e",
          6977 => x"af",
          6978 => x"ec",
          6979 => x"67",
          6980 => x"2e",
          6981 => x"82",
          6982 => x"8b",
          6983 => x"75",
          6984 => x"80",
          6985 => x"81",
          6986 => x"2e",
          6987 => x"80",
          6988 => x"38",
          6989 => x"0a",
          6990 => x"ff",
          6991 => x"55",
          6992 => x"86",
          6993 => x"8a",
          6994 => x"89",
          6995 => x"2a",
          6996 => x"77",
          6997 => x"59",
          6998 => x"81",
          6999 => x"81",
          7000 => x"25",
          7001 => x"55",
          7002 => x"8a",
          7003 => x"3d",
          7004 => x"81",
          7005 => x"ff",
          7006 => x"81",
          7007 => x"ec",
          7008 => x"38",
          7009 => x"70",
          7010 => x"85",
          7011 => x"56",
          7012 => x"38",
          7013 => x"55",
          7014 => x"75",
          7015 => x"38",
          7016 => x"70",
          7017 => x"ff",
          7018 => x"8c",
          7019 => x"78",
          7020 => x"8a",
          7021 => x"81",
          7022 => x"06",
          7023 => x"80",
          7024 => x"77",
          7025 => x"74",
          7026 => x"94",
          7027 => x"06",
          7028 => x"2e",
          7029 => x"77",
          7030 => x"93",
          7031 => x"74",
          7032 => x"d4",
          7033 => x"7d",
          7034 => x"81",
          7035 => x"38",
          7036 => x"66",
          7037 => x"81",
          7038 => x"d8",
          7039 => x"74",
          7040 => x"38",
          7041 => x"98",
          7042 => x"d8",
          7043 => x"82",
          7044 => x"57",
          7045 => x"80",
          7046 => x"76",
          7047 => x"38",
          7048 => x"51",
          7049 => x"3f",
          7050 => x"08",
          7051 => x"87",
          7052 => x"5e",
          7053 => x"80",
          7054 => x"ec",
          7055 => x"8a",
          7056 => x"fd",
          7057 => x"75",
          7058 => x"38",
          7059 => x"78",
          7060 => x"8c",
          7061 => x"0b",
          7062 => x"22",
          7063 => x"80",
          7064 => x"74",
          7065 => x"38",
          7066 => x"56",
          7067 => x"17",
          7068 => x"57",
          7069 => x"2e",
          7070 => x"75",
          7071 => x"79",
          7072 => x"fe",
          7073 => x"82",
          7074 => x"82",
          7075 => x"05",
          7076 => x"82",
          7077 => x"9f",
          7078 => x"38",
          7079 => x"85",
          7080 => x"2b",
          7081 => x"08",
          7082 => x"73",
          7083 => x"5a",
          7084 => x"83",
          7085 => x"2a",
          7086 => x"a0",
          7087 => x"7d",
          7088 => x"69",
          7089 => x"05",
          7090 => x"05",
          7091 => x"74",
          7092 => x"59",
          7093 => x"7d",
          7094 => x"81",
          7095 => x"76",
          7096 => x"41",
          7097 => x"76",
          7098 => x"84",
          7099 => x"62",
          7100 => x"51",
          7101 => x"26",
          7102 => x"75",
          7103 => x"31",
          7104 => x"65",
          7105 => x"fe",
          7106 => x"82",
          7107 => x"58",
          7108 => x"09",
          7109 => x"38",
          7110 => x"08",
          7111 => x"26",
          7112 => x"78",
          7113 => x"79",
          7114 => x"78",
          7115 => x"86",
          7116 => x"82",
          7117 => x"06",
          7118 => x"83",
          7119 => x"82",
          7120 => x"27",
          7121 => x"8f",
          7122 => x"55",
          7123 => x"26",
          7124 => x"59",
          7125 => x"62",
          7126 => x"74",
          7127 => x"38",
          7128 => x"81",
          7129 => x"ec",
          7130 => x"26",
          7131 => x"86",
          7132 => x"1a",
          7133 => x"79",
          7134 => x"38",
          7135 => x"80",
          7136 => x"2e",
          7137 => x"83",
          7138 => x"9f",
          7139 => x"8b",
          7140 => x"06",
          7141 => x"74",
          7142 => x"84",
          7143 => x"52",
          7144 => x"a1",
          7145 => x"53",
          7146 => x"52",
          7147 => x"a1",
          7148 => x"80",
          7149 => x"51",
          7150 => x"3f",
          7151 => x"34",
          7152 => x"ff",
          7153 => x"1b",
          7154 => x"d8",
          7155 => x"90",
          7156 => x"83",
          7157 => x"81",
          7158 => x"2a",
          7159 => x"54",
          7160 => x"1b",
          7161 => x"bc",
          7162 => x"74",
          7163 => x"26",
          7164 => x"83",
          7165 => x"52",
          7166 => x"ff",
          7167 => x"8a",
          7168 => x"a0",
          7169 => x"a0",
          7170 => x"0b",
          7171 => x"bf",
          7172 => x"51",
          7173 => x"3f",
          7174 => x"9a",
          7175 => x"a0",
          7176 => x"52",
          7177 => x"ff",
          7178 => x"7d",
          7179 => x"81",
          7180 => x"38",
          7181 => x"0a",
          7182 => x"1b",
          7183 => x"82",
          7184 => x"a4",
          7185 => x"9f",
          7186 => x"52",
          7187 => x"ff",
          7188 => x"81",
          7189 => x"51",
          7190 => x"3f",
          7191 => x"1b",
          7192 => x"c0",
          7193 => x"0b",
          7194 => x"34",
          7195 => x"c2",
          7196 => x"53",
          7197 => x"52",
          7198 => x"51",
          7199 => x"88",
          7200 => x"a7",
          7201 => x"9f",
          7202 => x"83",
          7203 => x"52",
          7204 => x"ff",
          7205 => x"ff",
          7206 => x"1c",
          7207 => x"a6",
          7208 => x"53",
          7209 => x"52",
          7210 => x"ff",
          7211 => x"82",
          7212 => x"83",
          7213 => x"52",
          7214 => x"e8",
          7215 => x"60",
          7216 => x"7e",
          7217 => x"8b",
          7218 => x"82",
          7219 => x"83",
          7220 => x"83",
          7221 => x"06",
          7222 => x"75",
          7223 => x"05",
          7224 => x"7e",
          7225 => x"eb",
          7226 => x"53",
          7227 => x"51",
          7228 => x"3f",
          7229 => x"a4",
          7230 => x"51",
          7231 => x"3f",
          7232 => x"e4",
          7233 => x"e4",
          7234 => x"9e",
          7235 => x"18",
          7236 => x"1b",
          7237 => x"aa",
          7238 => x"83",
          7239 => x"ff",
          7240 => x"82",
          7241 => x"78",
          7242 => x"f8",
          7243 => x"60",
          7244 => x"7a",
          7245 => x"ff",
          7246 => x"75",
          7247 => x"53",
          7248 => x"51",
          7249 => x"3f",
          7250 => x"52",
          7251 => x"9e",
          7252 => x"56",
          7253 => x"83",
          7254 => x"06",
          7255 => x"52",
          7256 => x"9d",
          7257 => x"52",
          7258 => x"ff",
          7259 => x"f0",
          7260 => x"1b",
          7261 => x"87",
          7262 => x"55",
          7263 => x"83",
          7264 => x"74",
          7265 => x"ff",
          7266 => x"7c",
          7267 => x"74",
          7268 => x"38",
          7269 => x"54",
          7270 => x"52",
          7271 => x"99",
          7272 => x"85",
          7273 => x"87",
          7274 => x"53",
          7275 => x"08",
          7276 => x"ff",
          7277 => x"76",
          7278 => x"31",
          7279 => x"cd",
          7280 => x"58",
          7281 => x"ff",
          7282 => x"55",
          7283 => x"83",
          7284 => x"61",
          7285 => x"26",
          7286 => x"57",
          7287 => x"53",
          7288 => x"51",
          7289 => x"3f",
          7290 => x"08",
          7291 => x"76",
          7292 => x"31",
          7293 => x"db",
          7294 => x"7d",
          7295 => x"38",
          7296 => x"83",
          7297 => x"8a",
          7298 => x"7d",
          7299 => x"38",
          7300 => x"81",
          7301 => x"80",
          7302 => x"80",
          7303 => x"7a",
          7304 => x"f0",
          7305 => x"d5",
          7306 => x"ff",
          7307 => x"83",
          7308 => x"77",
          7309 => x"0b",
          7310 => x"81",
          7311 => x"34",
          7312 => x"34",
          7313 => x"34",
          7314 => x"56",
          7315 => x"52",
          7316 => x"b9",
          7317 => x"0b",
          7318 => x"82",
          7319 => x"82",
          7320 => x"56",
          7321 => x"34",
          7322 => x"08",
          7323 => x"60",
          7324 => x"1b",
          7325 => x"ca",
          7326 => x"83",
          7327 => x"ff",
          7328 => x"81",
          7329 => x"7a",
          7330 => x"ff",
          7331 => x"81",
          7332 => x"ec",
          7333 => x"80",
          7334 => x"7e",
          7335 => x"97",
          7336 => x"82",
          7337 => x"90",
          7338 => x"8e",
          7339 => x"81",
          7340 => x"82",
          7341 => x"56",
          7342 => x"ec",
          7343 => x"0d",
          7344 => x"0d",
          7345 => x"59",
          7346 => x"ff",
          7347 => x"57",
          7348 => x"b4",
          7349 => x"f8",
          7350 => x"81",
          7351 => x"52",
          7352 => x"c0",
          7353 => x"2e",
          7354 => x"9c",
          7355 => x"33",
          7356 => x"2e",
          7357 => x"76",
          7358 => x"58",
          7359 => x"57",
          7360 => x"09",
          7361 => x"38",
          7362 => x"78",
          7363 => x"38",
          7364 => x"82",
          7365 => x"8d",
          7366 => x"f7",
          7367 => x"02",
          7368 => x"05",
          7369 => x"77",
          7370 => x"81",
          7371 => x"8d",
          7372 => x"e7",
          7373 => x"08",
          7374 => x"24",
          7375 => x"88",
          7376 => x"17",
          7377 => x"59",
          7378 => x"81",
          7379 => x"76",
          7380 => x"8b",
          7381 => x"54",
          7382 => x"17",
          7383 => x"51",
          7384 => x"79",
          7385 => x"09",
          7386 => x"72",
          7387 => x"70",
          7388 => x"53",
          7389 => x"75",
          7390 => x"81",
          7391 => x"0c",
          7392 => x"04",
          7393 => x"79",
          7394 => x"56",
          7395 => x"24",
          7396 => x"3d",
          7397 => x"74",
          7398 => x"52",
          7399 => x"cb",
          7400 => x"85",
          7401 => x"38",
          7402 => x"78",
          7403 => x"06",
          7404 => x"16",
          7405 => x"39",
          7406 => x"82",
          7407 => x"89",
          7408 => x"fd",
          7409 => x"54",
          7410 => x"80",
          7411 => x"ff",
          7412 => x"76",
          7413 => x"3d",
          7414 => x"3d",
          7415 => x"e3",
          7416 => x"53",
          7417 => x"53",
          7418 => x"3f",
          7419 => x"51",
          7420 => x"72",
          7421 => x"3f",
          7422 => x"04",
          7423 => x"ff",
          7424 => x"ff",
          7425 => x"00",
          7426 => x"ff",
          7427 => x"11",
          7428 => x"11",
          7429 => x"11",
          7430 => x"11",
          7431 => x"11",
          7432 => x"11",
          7433 => x"11",
          7434 => x"11",
          7435 => x"11",
          7436 => x"11",
          7437 => x"11",
          7438 => x"11",
          7439 => x"11",
          7440 => x"11",
          7441 => x"11",
          7442 => x"11",
          7443 => x"11",
          7444 => x"11",
          7445 => x"11",
          7446 => x"11",
          7447 => x"26",
          7448 => x"26",
          7449 => x"26",
          7450 => x"26",
          7451 => x"26",
          7452 => x"32",
          7453 => x"33",
          7454 => x"34",
          7455 => x"36",
          7456 => x"33",
          7457 => x"31",
          7458 => x"35",
          7459 => x"36",
          7460 => x"35",
          7461 => x"36",
          7462 => x"35",
          7463 => x"34",
          7464 => x"31",
          7465 => x"34",
          7466 => x"34",
          7467 => x"35",
          7468 => x"31",
          7469 => x"31",
          7470 => x"35",
          7471 => x"36",
          7472 => x"36",
          7473 => x"36",
          7474 => x"6e",
          7475 => x"00",
          7476 => x"6f",
          7477 => x"00",
          7478 => x"6e",
          7479 => x"00",
          7480 => x"6f",
          7481 => x"00",
          7482 => x"78",
          7483 => x"00",
          7484 => x"6c",
          7485 => x"00",
          7486 => x"6f",
          7487 => x"00",
          7488 => x"69",
          7489 => x"00",
          7490 => x"75",
          7491 => x"00",
          7492 => x"62",
          7493 => x"68",
          7494 => x"77",
          7495 => x"64",
          7496 => x"65",
          7497 => x"64",
          7498 => x"65",
          7499 => x"6c",
          7500 => x"00",
          7501 => x"70",
          7502 => x"73",
          7503 => x"74",
          7504 => x"73",
          7505 => x"00",
          7506 => x"66",
          7507 => x"00",
          7508 => x"73",
          7509 => x"00",
          7510 => x"61",
          7511 => x"00",
          7512 => x"61",
          7513 => x"00",
          7514 => x"6c",
          7515 => x"00",
          7516 => x"00",
          7517 => x"73",
          7518 => x"72",
          7519 => x"0a",
          7520 => x"74",
          7521 => x"61",
          7522 => x"72",
          7523 => x"2e",
          7524 => x"00",
          7525 => x"73",
          7526 => x"6f",
          7527 => x"65",
          7528 => x"2e",
          7529 => x"00",
          7530 => x"20",
          7531 => x"65",
          7532 => x"75",
          7533 => x"0a",
          7534 => x"20",
          7535 => x"68",
          7536 => x"75",
          7537 => x"0a",
          7538 => x"76",
          7539 => x"64",
          7540 => x"6c",
          7541 => x"6d",
          7542 => x"00",
          7543 => x"63",
          7544 => x"20",
          7545 => x"69",
          7546 => x"0a",
          7547 => x"6c",
          7548 => x"6c",
          7549 => x"64",
          7550 => x"78",
          7551 => x"73",
          7552 => x"00",
          7553 => x"6c",
          7554 => x"61",
          7555 => x"65",
          7556 => x"76",
          7557 => x"64",
          7558 => x"00",
          7559 => x"20",
          7560 => x"77",
          7561 => x"65",
          7562 => x"6f",
          7563 => x"74",
          7564 => x"0a",
          7565 => x"69",
          7566 => x"6e",
          7567 => x"65",
          7568 => x"73",
          7569 => x"76",
          7570 => x"64",
          7571 => x"00",
          7572 => x"73",
          7573 => x"6f",
          7574 => x"6e",
          7575 => x"65",
          7576 => x"00",
          7577 => x"20",
          7578 => x"70",
          7579 => x"62",
          7580 => x"66",
          7581 => x"73",
          7582 => x"65",
          7583 => x"6f",
          7584 => x"20",
          7585 => x"64",
          7586 => x"2e",
          7587 => x"00",
          7588 => x"72",
          7589 => x"20",
          7590 => x"72",
          7591 => x"2e",
          7592 => x"00",
          7593 => x"6d",
          7594 => x"74",
          7595 => x"70",
          7596 => x"74",
          7597 => x"20",
          7598 => x"63",
          7599 => x"65",
          7600 => x"00",
          7601 => x"6c",
          7602 => x"73",
          7603 => x"63",
          7604 => x"2e",
          7605 => x"00",
          7606 => x"73",
          7607 => x"69",
          7608 => x"6e",
          7609 => x"65",
          7610 => x"79",
          7611 => x"00",
          7612 => x"6f",
          7613 => x"6e",
          7614 => x"70",
          7615 => x"66",
          7616 => x"73",
          7617 => x"00",
          7618 => x"72",
          7619 => x"74",
          7620 => x"20",
          7621 => x"6f",
          7622 => x"63",
          7623 => x"00",
          7624 => x"63",
          7625 => x"73",
          7626 => x"00",
          7627 => x"6b",
          7628 => x"6e",
          7629 => x"72",
          7630 => x"0a",
          7631 => x"6c",
          7632 => x"79",
          7633 => x"20",
          7634 => x"61",
          7635 => x"6c",
          7636 => x"79",
          7637 => x"2f",
          7638 => x"2e",
          7639 => x"00",
          7640 => x"61",
          7641 => x"00",
          7642 => x"38",
          7643 => x"00",
          7644 => x"20",
          7645 => x"34",
          7646 => x"00",
          7647 => x"20",
          7648 => x"20",
          7649 => x"00",
          7650 => x"32",
          7651 => x"00",
          7652 => x"00",
          7653 => x"00",
          7654 => x"0a",
          7655 => x"53",
          7656 => x"2a",
          7657 => x"20",
          7658 => x"00",
          7659 => x"2f",
          7660 => x"32",
          7661 => x"00",
          7662 => x"2e",
          7663 => x"00",
          7664 => x"50",
          7665 => x"72",
          7666 => x"25",
          7667 => x"29",
          7668 => x"20",
          7669 => x"2a",
          7670 => x"00",
          7671 => x"55",
          7672 => x"74",
          7673 => x"75",
          7674 => x"48",
          7675 => x"6c",
          7676 => x"00",
          7677 => x"6d",
          7678 => x"69",
          7679 => x"72",
          7680 => x"74",
          7681 => x"00",
          7682 => x"32",
          7683 => x"74",
          7684 => x"75",
          7685 => x"00",
          7686 => x"43",
          7687 => x"52",
          7688 => x"6e",
          7689 => x"72",
          7690 => x"0a",
          7691 => x"43",
          7692 => x"57",
          7693 => x"6e",
          7694 => x"72",
          7695 => x"0a",
          7696 => x"52",
          7697 => x"52",
          7698 => x"6e",
          7699 => x"72",
          7700 => x"0a",
          7701 => x"52",
          7702 => x"54",
          7703 => x"6e",
          7704 => x"72",
          7705 => x"0a",
          7706 => x"52",
          7707 => x"52",
          7708 => x"6e",
          7709 => x"72",
          7710 => x"0a",
          7711 => x"52",
          7712 => x"54",
          7713 => x"6e",
          7714 => x"72",
          7715 => x"0a",
          7716 => x"74",
          7717 => x"67",
          7718 => x"20",
          7719 => x"65",
          7720 => x"2e",
          7721 => x"00",
          7722 => x"61",
          7723 => x"6e",
          7724 => x"69",
          7725 => x"2e",
          7726 => x"00",
          7727 => x"74",
          7728 => x"65",
          7729 => x"61",
          7730 => x"00",
          7731 => x"53",
          7732 => x"74",
          7733 => x"00",
          7734 => x"69",
          7735 => x"20",
          7736 => x"69",
          7737 => x"69",
          7738 => x"73",
          7739 => x"64",
          7740 => x"72",
          7741 => x"2c",
          7742 => x"65",
          7743 => x"20",
          7744 => x"74",
          7745 => x"6e",
          7746 => x"6c",
          7747 => x"00",
          7748 => x"00",
          7749 => x"65",
          7750 => x"6e",
          7751 => x"2e",
          7752 => x"00",
          7753 => x"70",
          7754 => x"67",
          7755 => x"00",
          7756 => x"6d",
          7757 => x"69",
          7758 => x"2e",
          7759 => x"00",
          7760 => x"38",
          7761 => x"25",
          7762 => x"29",
          7763 => x"30",
          7764 => x"28",
          7765 => x"78",
          7766 => x"00",
          7767 => x"6d",
          7768 => x"65",
          7769 => x"79",
          7770 => x"00",
          7771 => x"6f",
          7772 => x"65",
          7773 => x"0a",
          7774 => x"38",
          7775 => x"30",
          7776 => x"00",
          7777 => x"3f",
          7778 => x"00",
          7779 => x"38",
          7780 => x"30",
          7781 => x"00",
          7782 => x"38",
          7783 => x"30",
          7784 => x"00",
          7785 => x"65",
          7786 => x"69",
          7787 => x"63",
          7788 => x"20",
          7789 => x"30",
          7790 => x"2e",
          7791 => x"00",
          7792 => x"6c",
          7793 => x"67",
          7794 => x"64",
          7795 => x"20",
          7796 => x"78",
          7797 => x"2e",
          7798 => x"00",
          7799 => x"6c",
          7800 => x"65",
          7801 => x"6e",
          7802 => x"63",
          7803 => x"20",
          7804 => x"29",
          7805 => x"00",
          7806 => x"73",
          7807 => x"74",
          7808 => x"20",
          7809 => x"6c",
          7810 => x"74",
          7811 => x"2e",
          7812 => x"00",
          7813 => x"6c",
          7814 => x"65",
          7815 => x"74",
          7816 => x"2e",
          7817 => x"00",
          7818 => x"55",
          7819 => x"6e",
          7820 => x"3a",
          7821 => x"5c",
          7822 => x"25",
          7823 => x"00",
          7824 => x"3a",
          7825 => x"5c",
          7826 => x"00",
          7827 => x"3a",
          7828 => x"00",
          7829 => x"64",
          7830 => x"6d",
          7831 => x"64",
          7832 => x"00",
          7833 => x"6e",
          7834 => x"67",
          7835 => x"0a",
          7836 => x"61",
          7837 => x"6e",
          7838 => x"6e",
          7839 => x"72",
          7840 => x"73",
          7841 => x"0a",
          7842 => x"2f",
          7843 => x"25",
          7844 => x"64",
          7845 => x"3a",
          7846 => x"25",
          7847 => x"0a",
          7848 => x"43",
          7849 => x"6e",
          7850 => x"75",
          7851 => x"69",
          7852 => x"00",
          7853 => x"66",
          7854 => x"20",
          7855 => x"20",
          7856 => x"66",
          7857 => x"00",
          7858 => x"44",
          7859 => x"63",
          7860 => x"69",
          7861 => x"65",
          7862 => x"74",
          7863 => x"0a",
          7864 => x"20",
          7865 => x"20",
          7866 => x"41",
          7867 => x"28",
          7868 => x"58",
          7869 => x"38",
          7870 => x"0a",
          7871 => x"20",
          7872 => x"52",
          7873 => x"20",
          7874 => x"28",
          7875 => x"58",
          7876 => x"38",
          7877 => x"0a",
          7878 => x"20",
          7879 => x"53",
          7880 => x"52",
          7881 => x"28",
          7882 => x"58",
          7883 => x"38",
          7884 => x"0a",
          7885 => x"20",
          7886 => x"41",
          7887 => x"20",
          7888 => x"28",
          7889 => x"58",
          7890 => x"38",
          7891 => x"0a",
          7892 => x"20",
          7893 => x"4d",
          7894 => x"20",
          7895 => x"28",
          7896 => x"58",
          7897 => x"38",
          7898 => x"0a",
          7899 => x"20",
          7900 => x"20",
          7901 => x"44",
          7902 => x"28",
          7903 => x"69",
          7904 => x"20",
          7905 => x"32",
          7906 => x"0a",
          7907 => x"20",
          7908 => x"4d",
          7909 => x"20",
          7910 => x"28",
          7911 => x"65",
          7912 => x"20",
          7913 => x"32",
          7914 => x"0a",
          7915 => x"20",
          7916 => x"54",
          7917 => x"54",
          7918 => x"28",
          7919 => x"6e",
          7920 => x"73",
          7921 => x"32",
          7922 => x"0a",
          7923 => x"20",
          7924 => x"53",
          7925 => x"4e",
          7926 => x"55",
          7927 => x"00",
          7928 => x"20",
          7929 => x"20",
          7930 => x"0a",
          7931 => x"20",
          7932 => x"43",
          7933 => x"00",
          7934 => x"20",
          7935 => x"32",
          7936 => x"00",
          7937 => x"20",
          7938 => x"49",
          7939 => x"00",
          7940 => x"64",
          7941 => x"73",
          7942 => x"0a",
          7943 => x"20",
          7944 => x"55",
          7945 => x"73",
          7946 => x"56",
          7947 => x"6f",
          7948 => x"64",
          7949 => x"73",
          7950 => x"20",
          7951 => x"58",
          7952 => x"00",
          7953 => x"20",
          7954 => x"55",
          7955 => x"6d",
          7956 => x"20",
          7957 => x"72",
          7958 => x"64",
          7959 => x"73",
          7960 => x"20",
          7961 => x"58",
          7962 => x"00",
          7963 => x"20",
          7964 => x"61",
          7965 => x"53",
          7966 => x"74",
          7967 => x"64",
          7968 => x"73",
          7969 => x"20",
          7970 => x"20",
          7971 => x"58",
          7972 => x"00",
          7973 => x"73",
          7974 => x"00",
          7975 => x"20",
          7976 => x"55",
          7977 => x"20",
          7978 => x"20",
          7979 => x"20",
          7980 => x"20",
          7981 => x"20",
          7982 => x"20",
          7983 => x"58",
          7984 => x"00",
          7985 => x"20",
          7986 => x"73",
          7987 => x"20",
          7988 => x"63",
          7989 => x"72",
          7990 => x"20",
          7991 => x"20",
          7992 => x"20",
          7993 => x"25",
          7994 => x"4d",
          7995 => x"00",
          7996 => x"20",
          7997 => x"52",
          7998 => x"43",
          7999 => x"6b",
          8000 => x"65",
          8001 => x"20",
          8002 => x"20",
          8003 => x"20",
          8004 => x"25",
          8005 => x"4d",
          8006 => x"00",
          8007 => x"20",
          8008 => x"73",
          8009 => x"6e",
          8010 => x"44",
          8011 => x"20",
          8012 => x"63",
          8013 => x"72",
          8014 => x"20",
          8015 => x"25",
          8016 => x"4d",
          8017 => x"00",
          8018 => x"61",
          8019 => x"00",
          8020 => x"64",
          8021 => x"00",
          8022 => x"65",
          8023 => x"00",
          8024 => x"4f",
          8025 => x"4f",
          8026 => x"00",
          8027 => x"6b",
          8028 => x"6e",
          8029 => x"7e",
          8030 => x"00",
          8031 => x"00",
          8032 => x"7e",
          8033 => x"00",
          8034 => x"00",
          8035 => x"7e",
          8036 => x"00",
          8037 => x"00",
          8038 => x"7e",
          8039 => x"00",
          8040 => x"00",
          8041 => x"7e",
          8042 => x"00",
          8043 => x"00",
          8044 => x"7e",
          8045 => x"00",
          8046 => x"00",
          8047 => x"7e",
          8048 => x"00",
          8049 => x"00",
          8050 => x"7e",
          8051 => x"00",
          8052 => x"00",
          8053 => x"7e",
          8054 => x"00",
          8055 => x"00",
          8056 => x"7e",
          8057 => x"00",
          8058 => x"00",
          8059 => x"7e",
          8060 => x"00",
          8061 => x"00",
          8062 => x"7e",
          8063 => x"00",
          8064 => x"00",
          8065 => x"7e",
          8066 => x"00",
          8067 => x"00",
          8068 => x"7e",
          8069 => x"00",
          8070 => x"00",
          8071 => x"7e",
          8072 => x"00",
          8073 => x"00",
          8074 => x"7e",
          8075 => x"00",
          8076 => x"00",
          8077 => x"7e",
          8078 => x"00",
          8079 => x"00",
          8080 => x"7e",
          8081 => x"00",
          8082 => x"00",
          8083 => x"7e",
          8084 => x"00",
          8085 => x"00",
          8086 => x"7e",
          8087 => x"00",
          8088 => x"00",
          8089 => x"7e",
          8090 => x"00",
          8091 => x"00",
          8092 => x"7e",
          8093 => x"00",
          8094 => x"00",
          8095 => x"44",
          8096 => x"43",
          8097 => x"42",
          8098 => x"41",
          8099 => x"36",
          8100 => x"35",
          8101 => x"34",
          8102 => x"46",
          8103 => x"33",
          8104 => x"32",
          8105 => x"31",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"73",
          8118 => x"79",
          8119 => x"73",
          8120 => x"00",
          8121 => x"00",
          8122 => x"34",
          8123 => x"25",
          8124 => x"00",
          8125 => x"69",
          8126 => x"20",
          8127 => x"72",
          8128 => x"74",
          8129 => x"65",
          8130 => x"73",
          8131 => x"79",
          8132 => x"6c",
          8133 => x"6f",
          8134 => x"46",
          8135 => x"00",
          8136 => x"6e",
          8137 => x"20",
          8138 => x"6e",
          8139 => x"65",
          8140 => x"20",
          8141 => x"74",
          8142 => x"20",
          8143 => x"65",
          8144 => x"69",
          8145 => x"6c",
          8146 => x"2e",
          8147 => x"00",
          8148 => x"00",
          8149 => x"2b",
          8150 => x"3c",
          8151 => x"5b",
          8152 => x"00",
          8153 => x"54",
          8154 => x"54",
          8155 => x"00",
          8156 => x"90",
          8157 => x"4f",
          8158 => x"30",
          8159 => x"20",
          8160 => x"45",
          8161 => x"20",
          8162 => x"33",
          8163 => x"20",
          8164 => x"20",
          8165 => x"45",
          8166 => x"20",
          8167 => x"20",
          8168 => x"20",
          8169 => x"7f",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"45",
          8174 => x"8f",
          8175 => x"45",
          8176 => x"8e",
          8177 => x"92",
          8178 => x"55",
          8179 => x"9a",
          8180 => x"9e",
          8181 => x"4f",
          8182 => x"a6",
          8183 => x"aa",
          8184 => x"ae",
          8185 => x"b2",
          8186 => x"b6",
          8187 => x"ba",
          8188 => x"be",
          8189 => x"c2",
          8190 => x"c6",
          8191 => x"ca",
          8192 => x"ce",
          8193 => x"d2",
          8194 => x"d6",
          8195 => x"da",
          8196 => x"de",
          8197 => x"e2",
          8198 => x"e6",
          8199 => x"ea",
          8200 => x"ee",
          8201 => x"f2",
          8202 => x"f6",
          8203 => x"fa",
          8204 => x"fe",
          8205 => x"2c",
          8206 => x"5d",
          8207 => x"2a",
          8208 => x"3f",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"02",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"74",
          8220 => x"01",
          8221 => x"00",
          8222 => x"00",
          8223 => x"74",
          8224 => x"01",
          8225 => x"00",
          8226 => x"00",
          8227 => x"74",
          8228 => x"03",
          8229 => x"00",
          8230 => x"00",
          8231 => x"74",
          8232 => x"03",
          8233 => x"00",
          8234 => x"00",
          8235 => x"74",
          8236 => x"03",
          8237 => x"00",
          8238 => x"00",
          8239 => x"74",
          8240 => x"04",
          8241 => x"00",
          8242 => x"00",
          8243 => x"74",
          8244 => x"04",
          8245 => x"00",
          8246 => x"00",
          8247 => x"75",
          8248 => x"04",
          8249 => x"00",
          8250 => x"00",
          8251 => x"75",
          8252 => x"04",
          8253 => x"00",
          8254 => x"00",
          8255 => x"75",
          8256 => x"04",
          8257 => x"00",
          8258 => x"00",
          8259 => x"75",
          8260 => x"04",
          8261 => x"00",
          8262 => x"00",
          8263 => x"75",
          8264 => x"04",
          8265 => x"00",
          8266 => x"00",
          8267 => x"75",
          8268 => x"05",
          8269 => x"00",
          8270 => x"00",
          8271 => x"75",
          8272 => x"05",
          8273 => x"00",
          8274 => x"00",
          8275 => x"75",
          8276 => x"05",
          8277 => x"00",
          8278 => x"00",
          8279 => x"75",
          8280 => x"05",
          8281 => x"00",
          8282 => x"00",
          8283 => x"75",
          8284 => x"07",
          8285 => x"00",
          8286 => x"00",
          8287 => x"75",
          8288 => x"07",
          8289 => x"00",
          8290 => x"00",
          8291 => x"75",
          8292 => x"08",
          8293 => x"00",
          8294 => x"00",
          8295 => x"75",
          8296 => x"08",
          8297 => x"00",
          8298 => x"00",
          8299 => x"75",
          8300 => x"08",
          8301 => x"00",
          8302 => x"00",
          8303 => x"75",
          8304 => x"08",
          8305 => x"00",
          8306 => x"00",
          8307 => x"75",
          8308 => x"09",
          8309 => x"00",
          8310 => x"00",
          8311 => x"75",
          8312 => x"09",
          8313 => x"00",
          8314 => x"00",
          8315 => x"75",
          8316 => x"09",
          8317 => x"00",
          8318 => x"00",
          8319 => x"75",
          8320 => x"09",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"7f",
          8326 => x"00",
          8327 => x"7f",
          8328 => x"00",
          8329 => x"7f",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"ff",
          8334 => x"00",
          8335 => x"00",
          8336 => x"78",
          8337 => x"00",
          8338 => x"e1",
          8339 => x"e1",
          8340 => x"e1",
          8341 => x"00",
          8342 => x"01",
          8343 => x"01",
          8344 => x"10",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"7e",
          8371 => x"00",
          8372 => x"7e",
          8373 => x"00",
          8374 => x"7e",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"e7",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8e",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8f",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"90",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"91",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"92",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"82",
           389 => x"82",
           390 => x"80",
           391 => x"82",
           392 => x"82",
           393 => x"82",
           394 => x"80",
           395 => x"82",
           396 => x"82",
           397 => x"82",
           398 => x"80",
           399 => x"82",
           400 => x"82",
           401 => x"82",
           402 => x"80",
           403 => x"82",
           404 => x"82",
           405 => x"82",
           406 => x"80",
           407 => x"82",
           408 => x"82",
           409 => x"82",
           410 => x"80",
           411 => x"82",
           412 => x"82",
           413 => x"82",
           414 => x"80",
           415 => x"82",
           416 => x"82",
           417 => x"82",
           418 => x"80",
           419 => x"82",
           420 => x"82",
           421 => x"82",
           422 => x"80",
           423 => x"82",
           424 => x"82",
           425 => x"82",
           426 => x"80",
           427 => x"82",
           428 => x"82",
           429 => x"82",
           430 => x"80",
           431 => x"82",
           432 => x"82",
           433 => x"82",
           434 => x"80",
           435 => x"82",
           436 => x"82",
           437 => x"82",
           438 => x"80",
           439 => x"82",
           440 => x"82",
           441 => x"82",
           442 => x"80",
           443 => x"82",
           444 => x"82",
           445 => x"82",
           446 => x"bb",
           447 => x"85",
           448 => x"a0",
           449 => x"85",
           450 => x"bd",
           451 => x"f8",
           452 => x"90",
           453 => x"f8",
           454 => x"2d",
           455 => x"08",
           456 => x"04",
           457 => x"0c",
           458 => x"2d",
           459 => x"08",
           460 => x"04",
           461 => x"0c",
           462 => x"2d",
           463 => x"08",
           464 => x"04",
           465 => x"0c",
           466 => x"2d",
           467 => x"08",
           468 => x"04",
           469 => x"0c",
           470 => x"2d",
           471 => x"08",
           472 => x"04",
           473 => x"0c",
           474 => x"2d",
           475 => x"08",
           476 => x"04",
           477 => x"0c",
           478 => x"2d",
           479 => x"08",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"04",
           497 => x"0c",
           498 => x"2d",
           499 => x"08",
           500 => x"04",
           501 => x"0c",
           502 => x"2d",
           503 => x"08",
           504 => x"04",
           505 => x"0c",
           506 => x"2d",
           507 => x"08",
           508 => x"04",
           509 => x"0c",
           510 => x"2d",
           511 => x"08",
           512 => x"04",
           513 => x"0c",
           514 => x"2d",
           515 => x"08",
           516 => x"04",
           517 => x"0c",
           518 => x"2d",
           519 => x"08",
           520 => x"04",
           521 => x"0c",
           522 => x"2d",
           523 => x"08",
           524 => x"04",
           525 => x"0c",
           526 => x"2d",
           527 => x"08",
           528 => x"04",
           529 => x"0c",
           530 => x"2d",
           531 => x"08",
           532 => x"04",
           533 => x"0c",
           534 => x"2d",
           535 => x"08",
           536 => x"04",
           537 => x"0c",
           538 => x"2d",
           539 => x"08",
           540 => x"04",
           541 => x"0c",
           542 => x"2d",
           543 => x"08",
           544 => x"04",
           545 => x"0c",
           546 => x"2d",
           547 => x"08",
           548 => x"04",
           549 => x"0c",
           550 => x"2d",
           551 => x"08",
           552 => x"04",
           553 => x"0c",
           554 => x"2d",
           555 => x"08",
           556 => x"04",
           557 => x"0c",
           558 => x"2d",
           559 => x"08",
           560 => x"04",
           561 => x"0c",
           562 => x"2d",
           563 => x"08",
           564 => x"04",
           565 => x"0c",
           566 => x"2d",
           567 => x"08",
           568 => x"04",
           569 => x"0c",
           570 => x"2d",
           571 => x"08",
           572 => x"04",
           573 => x"0c",
           574 => x"2d",
           575 => x"08",
           576 => x"04",
           577 => x"0c",
           578 => x"82",
           579 => x"82",
           580 => x"82",
           581 => x"bd",
           582 => x"85",
           583 => x"a0",
           584 => x"85",
           585 => x"c0",
           586 => x"85",
           587 => x"a0",
           588 => x"85",
           589 => x"fd",
           590 => x"f8",
           591 => x"90",
           592 => x"00",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"10",
           598 => x"10",
           599 => x"10",
           600 => x"10",
           601 => x"00",
           602 => x"ff",
           603 => x"06",
           604 => x"83",
           605 => x"10",
           606 => x"fc",
           607 => x"51",
           608 => x"80",
           609 => x"ff",
           610 => x"06",
           611 => x"52",
           612 => x"0a",
           613 => x"38",
           614 => x"51",
           615 => x"ec",
           616 => x"a8",
           617 => x"80",
           618 => x"05",
           619 => x"0b",
           620 => x"04",
           621 => x"ba",
           622 => x"82",
           623 => x"02",
           624 => x"0c",
           625 => x"82",
           626 => x"88",
           627 => x"85",
           628 => x"05",
           629 => x"f8",
           630 => x"08",
           631 => x"82",
           632 => x"fc",
           633 => x"05",
           634 => x"08",
           635 => x"70",
           636 => x"51",
           637 => x"2e",
           638 => x"39",
           639 => x"08",
           640 => x"ff",
           641 => x"f8",
           642 => x"0c",
           643 => x"08",
           644 => x"82",
           645 => x"88",
           646 => x"70",
           647 => x"0c",
           648 => x"0d",
           649 => x"0c",
           650 => x"f8",
           651 => x"85",
           652 => x"3d",
           653 => x"f8",
           654 => x"08",
           655 => x"08",
           656 => x"82",
           657 => x"8c",
           658 => x"71",
           659 => x"f8",
           660 => x"08",
           661 => x"85",
           662 => x"05",
           663 => x"f8",
           664 => x"08",
           665 => x"72",
           666 => x"f8",
           667 => x"08",
           668 => x"85",
           669 => x"05",
           670 => x"ff",
           671 => x"80",
           672 => x"ff",
           673 => x"85",
           674 => x"05",
           675 => x"85",
           676 => x"84",
           677 => x"85",
           678 => x"82",
           679 => x"02",
           680 => x"0c",
           681 => x"82",
           682 => x"88",
           683 => x"85",
           684 => x"05",
           685 => x"f8",
           686 => x"08",
           687 => x"08",
           688 => x"82",
           689 => x"90",
           690 => x"2e",
           691 => x"82",
           692 => x"90",
           693 => x"05",
           694 => x"08",
           695 => x"82",
           696 => x"90",
           697 => x"05",
           698 => x"08",
           699 => x"82",
           700 => x"90",
           701 => x"2e",
           702 => x"85",
           703 => x"05",
           704 => x"33",
           705 => x"08",
           706 => x"81",
           707 => x"f8",
           708 => x"0c",
           709 => x"08",
           710 => x"52",
           711 => x"34",
           712 => x"08",
           713 => x"81",
           714 => x"f8",
           715 => x"0c",
           716 => x"82",
           717 => x"88",
           718 => x"82",
           719 => x"51",
           720 => x"82",
           721 => x"04",
           722 => x"08",
           723 => x"f8",
           724 => x"0d",
           725 => x"08",
           726 => x"80",
           727 => x"38",
           728 => x"08",
           729 => x"52",
           730 => x"85",
           731 => x"05",
           732 => x"82",
           733 => x"8c",
           734 => x"85",
           735 => x"05",
           736 => x"72",
           737 => x"53",
           738 => x"71",
           739 => x"38",
           740 => x"82",
           741 => x"88",
           742 => x"71",
           743 => x"f8",
           744 => x"08",
           745 => x"85",
           746 => x"05",
           747 => x"ff",
           748 => x"70",
           749 => x"0b",
           750 => x"08",
           751 => x"81",
           752 => x"85",
           753 => x"05",
           754 => x"82",
           755 => x"90",
           756 => x"85",
           757 => x"05",
           758 => x"84",
           759 => x"39",
           760 => x"08",
           761 => x"80",
           762 => x"38",
           763 => x"08",
           764 => x"70",
           765 => x"70",
           766 => x"0b",
           767 => x"08",
           768 => x"80",
           769 => x"85",
           770 => x"05",
           771 => x"82",
           772 => x"8c",
           773 => x"85",
           774 => x"05",
           775 => x"52",
           776 => x"38",
           777 => x"85",
           778 => x"05",
           779 => x"82",
           780 => x"88",
           781 => x"33",
           782 => x"08",
           783 => x"70",
           784 => x"31",
           785 => x"f8",
           786 => x"0c",
           787 => x"52",
           788 => x"80",
           789 => x"f8",
           790 => x"0c",
           791 => x"08",
           792 => x"82",
           793 => x"85",
           794 => x"85",
           795 => x"82",
           796 => x"02",
           797 => x"0c",
           798 => x"82",
           799 => x"88",
           800 => x"85",
           801 => x"05",
           802 => x"f8",
           803 => x"08",
           804 => x"d4",
           805 => x"f8",
           806 => x"08",
           807 => x"85",
           808 => x"05",
           809 => x"f8",
           810 => x"08",
           811 => x"85",
           812 => x"05",
           813 => x"f8",
           814 => x"08",
           815 => x"38",
           816 => x"08",
           817 => x"51",
           818 => x"f8",
           819 => x"08",
           820 => x"71",
           821 => x"f8",
           822 => x"08",
           823 => x"85",
           824 => x"05",
           825 => x"39",
           826 => x"08",
           827 => x"70",
           828 => x"0c",
           829 => x"0d",
           830 => x"0c",
           831 => x"f8",
           832 => x"85",
           833 => x"3d",
           834 => x"82",
           835 => x"fc",
           836 => x"85",
           837 => x"05",
           838 => x"b9",
           839 => x"f8",
           840 => x"08",
           841 => x"f8",
           842 => x"0c",
           843 => x"85",
           844 => x"05",
           845 => x"f8",
           846 => x"08",
           847 => x"0b",
           848 => x"08",
           849 => x"82",
           850 => x"f4",
           851 => x"85",
           852 => x"05",
           853 => x"f8",
           854 => x"08",
           855 => x"38",
           856 => x"08",
           857 => x"30",
           858 => x"08",
           859 => x"80",
           860 => x"f8",
           861 => x"0c",
           862 => x"08",
           863 => x"8a",
           864 => x"82",
           865 => x"f0",
           866 => x"85",
           867 => x"05",
           868 => x"f8",
           869 => x"0c",
           870 => x"85",
           871 => x"05",
           872 => x"85",
           873 => x"05",
           874 => x"c5",
           875 => x"ec",
           876 => x"85",
           877 => x"05",
           878 => x"85",
           879 => x"05",
           880 => x"90",
           881 => x"f8",
           882 => x"08",
           883 => x"f8",
           884 => x"0c",
           885 => x"08",
           886 => x"70",
           887 => x"0c",
           888 => x"0d",
           889 => x"0c",
           890 => x"f8",
           891 => x"85",
           892 => x"3d",
           893 => x"82",
           894 => x"fc",
           895 => x"85",
           896 => x"05",
           897 => x"99",
           898 => x"f8",
           899 => x"08",
           900 => x"f8",
           901 => x"0c",
           902 => x"85",
           903 => x"05",
           904 => x"f8",
           905 => x"08",
           906 => x"38",
           907 => x"08",
           908 => x"30",
           909 => x"08",
           910 => x"81",
           911 => x"f8",
           912 => x"08",
           913 => x"f8",
           914 => x"08",
           915 => x"3f",
           916 => x"08",
           917 => x"f8",
           918 => x"0c",
           919 => x"f8",
           920 => x"08",
           921 => x"38",
           922 => x"08",
           923 => x"30",
           924 => x"08",
           925 => x"82",
           926 => x"f8",
           927 => x"82",
           928 => x"54",
           929 => x"82",
           930 => x"04",
           931 => x"08",
           932 => x"f8",
           933 => x"0d",
           934 => x"85",
           935 => x"05",
           936 => x"f8",
           937 => x"08",
           938 => x"11",
           939 => x"82",
           940 => x"8c",
           941 => x"82",
           942 => x"fc",
           943 => x"82",
           944 => x"fc",
           945 => x"85",
           946 => x"05",
           947 => x"82",
           948 => x"88",
           949 => x"85",
           950 => x"05",
           951 => x"85",
           952 => x"05",
           953 => x"51",
           954 => x"f8",
           955 => x"08",
           956 => x"38",
           957 => x"82",
           958 => x"fc",
           959 => x"82",
           960 => x"51",
           961 => x"82",
           962 => x"04",
           963 => x"08",
           964 => x"f8",
           965 => x"0d",
           966 => x"85",
           967 => x"05",
           968 => x"85",
           969 => x"05",
           970 => x"c5",
           971 => x"ec",
           972 => x"85",
           973 => x"85",
           974 => x"85",
           975 => x"82",
           976 => x"02",
           977 => x"0c",
           978 => x"81",
           979 => x"f8",
           980 => x"08",
           981 => x"f8",
           982 => x"08",
           983 => x"82",
           984 => x"70",
           985 => x"0c",
           986 => x"0d",
           987 => x"0c",
           988 => x"f8",
           989 => x"85",
           990 => x"3d",
           991 => x"82",
           992 => x"fc",
           993 => x"0b",
           994 => x"08",
           995 => x"82",
           996 => x"8c",
           997 => x"85",
           998 => x"05",
           999 => x"38",
          1000 => x"08",
          1001 => x"80",
          1002 => x"80",
          1003 => x"f8",
          1004 => x"08",
          1005 => x"82",
          1006 => x"8c",
          1007 => x"82",
          1008 => x"8c",
          1009 => x"85",
          1010 => x"05",
          1011 => x"85",
          1012 => x"05",
          1013 => x"39",
          1014 => x"08",
          1015 => x"80",
          1016 => x"38",
          1017 => x"08",
          1018 => x"82",
          1019 => x"88",
          1020 => x"ad",
          1021 => x"f8",
          1022 => x"08",
          1023 => x"08",
          1024 => x"31",
          1025 => x"08",
          1026 => x"82",
          1027 => x"f8",
          1028 => x"85",
          1029 => x"05",
          1030 => x"85",
          1031 => x"05",
          1032 => x"f8",
          1033 => x"08",
          1034 => x"85",
          1035 => x"05",
          1036 => x"f8",
          1037 => x"08",
          1038 => x"85",
          1039 => x"05",
          1040 => x"39",
          1041 => x"08",
          1042 => x"80",
          1043 => x"82",
          1044 => x"88",
          1045 => x"82",
          1046 => x"f4",
          1047 => x"91",
          1048 => x"f8",
          1049 => x"08",
          1050 => x"f8",
          1051 => x"0c",
          1052 => x"f8",
          1053 => x"08",
          1054 => x"0c",
          1055 => x"82",
          1056 => x"04",
          1057 => x"79",
          1058 => x"56",
          1059 => x"80",
          1060 => x"38",
          1061 => x"08",
          1062 => x"3f",
          1063 => x"08",
          1064 => x"85",
          1065 => x"80",
          1066 => x"33",
          1067 => x"2e",
          1068 => x"86",
          1069 => x"55",
          1070 => x"57",
          1071 => x"82",
          1072 => x"70",
          1073 => x"f1",
          1074 => x"85",
          1075 => x"74",
          1076 => x"51",
          1077 => x"82",
          1078 => x"8b",
          1079 => x"33",
          1080 => x"2e",
          1081 => x"81",
          1082 => x"ff",
          1083 => x"99",
          1084 => x"38",
          1085 => x"82",
          1086 => x"89",
          1087 => x"ff",
          1088 => x"52",
          1089 => x"81",
          1090 => x"82",
          1091 => x"e8",
          1092 => x"04",
          1093 => x"51",
          1094 => x"81",
          1095 => x"80",
          1096 => x"eb",
          1097 => x"f2",
          1098 => x"a8",
          1099 => x"39",
          1100 => x"51",
          1101 => x"81",
          1102 => x"80",
          1103 => x"eb",
          1104 => x"d6",
          1105 => x"ec",
          1106 => x"39",
          1107 => x"51",
          1108 => x"81",
          1109 => x"80",
          1110 => x"ec",
          1111 => x"39",
          1112 => x"51",
          1113 => x"ec",
          1114 => x"39",
          1115 => x"51",
          1116 => x"ed",
          1117 => x"39",
          1118 => x"51",
          1119 => x"ed",
          1120 => x"39",
          1121 => x"51",
          1122 => x"ee",
          1123 => x"39",
          1124 => x"51",
          1125 => x"ee",
          1126 => x"d1",
          1127 => x"0d",
          1128 => x"0d",
          1129 => x"56",
          1130 => x"26",
          1131 => x"e8",
          1132 => x"f9",
          1133 => x"52",
          1134 => x"08",
          1135 => x"87",
          1136 => x"51",
          1137 => x"82",
          1138 => x"52",
          1139 => x"bc",
          1140 => x"ec",
          1141 => x"53",
          1142 => x"ee",
          1143 => x"fd",
          1144 => x"0d",
          1145 => x"0d",
          1146 => x"05",
          1147 => x"33",
          1148 => x"68",
          1149 => x"05",
          1150 => x"73",
          1151 => x"59",
          1152 => x"77",
          1153 => x"83",
          1154 => x"74",
          1155 => x"81",
          1156 => x"55",
          1157 => x"81",
          1158 => x"53",
          1159 => x"3d",
          1160 => x"81",
          1161 => x"82",
          1162 => x"57",
          1163 => x"08",
          1164 => x"85",
          1165 => x"c0",
          1166 => x"82",
          1167 => x"59",
          1168 => x"05",
          1169 => x"53",
          1170 => x"51",
          1171 => x"3f",
          1172 => x"08",
          1173 => x"ec",
          1174 => x"7a",
          1175 => x"2e",
          1176 => x"19",
          1177 => x"59",
          1178 => x"3d",
          1179 => x"81",
          1180 => x"76",
          1181 => x"70",
          1182 => x"25",
          1183 => x"05",
          1184 => x"72",
          1185 => x"51",
          1186 => x"2e",
          1187 => x"ee",
          1188 => x"c0",
          1189 => x"52",
          1190 => x"85",
          1191 => x"75",
          1192 => x"0c",
          1193 => x"04",
          1194 => x"7b",
          1195 => x"b3",
          1196 => x"58",
          1197 => x"53",
          1198 => x"51",
          1199 => x"82",
          1200 => x"a4",
          1201 => x"2e",
          1202 => x"81",
          1203 => x"98",
          1204 => x"7f",
          1205 => x"ec",
          1206 => x"7d",
          1207 => x"82",
          1208 => x"57",
          1209 => x"04",
          1210 => x"ec",
          1211 => x"0d",
          1212 => x"0d",
          1213 => x"02",
          1214 => x"cf",
          1215 => x"73",
          1216 => x"5f",
          1217 => x"5e",
          1218 => x"81",
          1219 => x"ae",
          1220 => x"ee",
          1221 => x"d5",
          1222 => x"74",
          1223 => x"f4",
          1224 => x"2e",
          1225 => x"a0",
          1226 => x"80",
          1227 => x"18",
          1228 => x"27",
          1229 => x"22",
          1230 => x"f4",
          1231 => x"3f",
          1232 => x"ef",
          1233 => x"a5",
          1234 => x"55",
          1235 => x"18",
          1236 => x"27",
          1237 => x"08",
          1238 => x"e8",
          1239 => x"3f",
          1240 => x"ee",
          1241 => x"85",
          1242 => x"55",
          1243 => x"18",
          1244 => x"27",
          1245 => x"33",
          1246 => x"88",
          1247 => x"3f",
          1248 => x"ef",
          1249 => x"e5",
          1250 => x"55",
          1251 => x"80",
          1252 => x"39",
          1253 => x"51",
          1254 => x"80",
          1255 => x"27",
          1256 => x"18",
          1257 => x"53",
          1258 => x"7a",
          1259 => x"81",
          1260 => x"9f",
          1261 => x"38",
          1262 => x"73",
          1263 => x"ff",
          1264 => x"72",
          1265 => x"38",
          1266 => x"26",
          1267 => x"51",
          1268 => x"51",
          1269 => x"81",
          1270 => x"39",
          1271 => x"51",
          1272 => x"78",
          1273 => x"5c",
          1274 => x"3f",
          1275 => x"08",
          1276 => x"98",
          1277 => x"76",
          1278 => x"81",
          1279 => x"9b",
          1280 => x"85",
          1281 => x"2b",
          1282 => x"70",
          1283 => x"09",
          1284 => x"9b",
          1285 => x"81",
          1286 => x"07",
          1287 => x"06",
          1288 => x"59",
          1289 => x"80",
          1290 => x"38",
          1291 => x"09",
          1292 => x"38",
          1293 => x"39",
          1294 => x"72",
          1295 => x"c9",
          1296 => x"72",
          1297 => x"0c",
          1298 => x"04",
          1299 => x"02",
          1300 => x"81",
          1301 => x"81",
          1302 => x"55",
          1303 => x"82",
          1304 => x"51",
          1305 => x"81",
          1306 => x"81",
          1307 => x"82",
          1308 => x"52",
          1309 => x"51",
          1310 => x"74",
          1311 => x"38",
          1312 => x"86",
          1313 => x"fe",
          1314 => x"c0",
          1315 => x"53",
          1316 => x"81",
          1317 => x"3f",
          1318 => x"51",
          1319 => x"80",
          1320 => x"3f",
          1321 => x"70",
          1322 => x"52",
          1323 => x"92",
          1324 => x"96",
          1325 => x"ef",
          1326 => x"c2",
          1327 => x"96",
          1328 => x"82",
          1329 => x"06",
          1330 => x"80",
          1331 => x"81",
          1332 => x"3f",
          1333 => x"51",
          1334 => x"80",
          1335 => x"3f",
          1336 => x"70",
          1337 => x"52",
          1338 => x"92",
          1339 => x"96",
          1340 => x"f0",
          1341 => x"86",
          1342 => x"96",
          1343 => x"84",
          1344 => x"06",
          1345 => x"80",
          1346 => x"81",
          1347 => x"3f",
          1348 => x"51",
          1349 => x"80",
          1350 => x"3f",
          1351 => x"70",
          1352 => x"52",
          1353 => x"92",
          1354 => x"95",
          1355 => x"f0",
          1356 => x"ca",
          1357 => x"95",
          1358 => x"86",
          1359 => x"06",
          1360 => x"80",
          1361 => x"81",
          1362 => x"3f",
          1363 => x"51",
          1364 => x"80",
          1365 => x"3f",
          1366 => x"70",
          1367 => x"52",
          1368 => x"92",
          1369 => x"95",
          1370 => x"f0",
          1371 => x"8e",
          1372 => x"95",
          1373 => x"88",
          1374 => x"06",
          1375 => x"80",
          1376 => x"81",
          1377 => x"3f",
          1378 => x"51",
          1379 => x"80",
          1380 => x"3f",
          1381 => x"84",
          1382 => x"fb",
          1383 => x"02",
          1384 => x"05",
          1385 => x"56",
          1386 => x"75",
          1387 => x"3f",
          1388 => x"80",
          1389 => x"73",
          1390 => x"53",
          1391 => x"52",
          1392 => x"51",
          1393 => x"3f",
          1394 => x"08",
          1395 => x"70",
          1396 => x"08",
          1397 => x"82",
          1398 => x"51",
          1399 => x"0b",
          1400 => x"34",
          1401 => x"80",
          1402 => x"73",
          1403 => x"81",
          1404 => x"82",
          1405 => x"74",
          1406 => x"81",
          1407 => x"82",
          1408 => x"80",
          1409 => x"82",
          1410 => x"51",
          1411 => x"91",
          1412 => x"cc",
          1413 => x"99",
          1414 => x"0b",
          1415 => x"e8",
          1416 => x"82",
          1417 => x"54",
          1418 => x"09",
          1419 => x"38",
          1420 => x"53",
          1421 => x"51",
          1422 => x"80",
          1423 => x"ec",
          1424 => x"0d",
          1425 => x"0d",
          1426 => x"82",
          1427 => x"5f",
          1428 => x"7c",
          1429 => x"93",
          1430 => x"ec",
          1431 => x"06",
          1432 => x"2e",
          1433 => x"a1",
          1434 => x"d4",
          1435 => x"70",
          1436 => x"ff",
          1437 => x"78",
          1438 => x"f8",
          1439 => x"dd",
          1440 => x"ec",
          1441 => x"88",
          1442 => x"d8",
          1443 => x"39",
          1444 => x"5d",
          1445 => x"51",
          1446 => x"96",
          1447 => x"5a",
          1448 => x"79",
          1449 => x"3f",
          1450 => x"84",
          1451 => x"d4",
          1452 => x"ec",
          1453 => x"70",
          1454 => x"59",
          1455 => x"2e",
          1456 => x"78",
          1457 => x"b2",
          1458 => x"2e",
          1459 => x"78",
          1460 => x"38",
          1461 => x"ff",
          1462 => x"bc",
          1463 => x"38",
          1464 => x"78",
          1465 => x"83",
          1466 => x"80",
          1467 => x"cd",
          1468 => x"2e",
          1469 => x"8a",
          1470 => x"80",
          1471 => x"c3",
          1472 => x"f9",
          1473 => x"78",
          1474 => x"87",
          1475 => x"80",
          1476 => x"8c",
          1477 => x"39",
          1478 => x"2e",
          1479 => x"78",
          1480 => x"8b",
          1481 => x"82",
          1482 => x"38",
          1483 => x"78",
          1484 => x"89",
          1485 => x"e5",
          1486 => x"ff",
          1487 => x"ff",
          1488 => x"a8",
          1489 => x"85",
          1490 => x"2e",
          1491 => x"b4",
          1492 => x"11",
          1493 => x"05",
          1494 => x"3f",
          1495 => x"08",
          1496 => x"b0",
          1497 => x"fe",
          1498 => x"ff",
          1499 => x"a7",
          1500 => x"85",
          1501 => x"38",
          1502 => x"08",
          1503 => x"94",
          1504 => x"3f",
          1505 => x"5a",
          1506 => x"81",
          1507 => x"59",
          1508 => x"84",
          1509 => x"7a",
          1510 => x"38",
          1511 => x"b4",
          1512 => x"11",
          1513 => x"05",
          1514 => x"3f",
          1515 => x"08",
          1516 => x"e0",
          1517 => x"fe",
          1518 => x"ff",
          1519 => x"a7",
          1520 => x"85",
          1521 => x"2e",
          1522 => x"b4",
          1523 => x"11",
          1524 => x"05",
          1525 => x"3f",
          1526 => x"08",
          1527 => x"b4",
          1528 => x"a4",
          1529 => x"3f",
          1530 => x"63",
          1531 => x"38",
          1532 => x"70",
          1533 => x"33",
          1534 => x"81",
          1535 => x"39",
          1536 => x"80",
          1537 => x"84",
          1538 => x"c9",
          1539 => x"ec",
          1540 => x"fc",
          1541 => x"3d",
          1542 => x"53",
          1543 => x"51",
          1544 => x"82",
          1545 => x"80",
          1546 => x"38",
          1547 => x"f8",
          1548 => x"84",
          1549 => x"9d",
          1550 => x"ec",
          1551 => x"fc",
          1552 => x"f2",
          1553 => x"a5",
          1554 => x"79",
          1555 => x"38",
          1556 => x"7b",
          1557 => x"5b",
          1558 => x"91",
          1559 => x"7a",
          1560 => x"53",
          1561 => x"f2",
          1562 => x"f1",
          1563 => x"62",
          1564 => x"5a",
          1565 => x"f2",
          1566 => x"bb",
          1567 => x"ff",
          1568 => x"ff",
          1569 => x"a5",
          1570 => x"85",
          1571 => x"df",
          1572 => x"d8",
          1573 => x"80",
          1574 => x"82",
          1575 => x"44",
          1576 => x"82",
          1577 => x"59",
          1578 => x"88",
          1579 => x"98",
          1580 => x"39",
          1581 => x"33",
          1582 => x"2e",
          1583 => x"84",
          1584 => x"ab",
          1585 => x"db",
          1586 => x"80",
          1587 => x"82",
          1588 => x"44",
          1589 => x"84",
          1590 => x"78",
          1591 => x"38",
          1592 => x"08",
          1593 => x"82",
          1594 => x"fc",
          1595 => x"b4",
          1596 => x"11",
          1597 => x"05",
          1598 => x"3f",
          1599 => x"08",
          1600 => x"82",
          1601 => x"59",
          1602 => x"89",
          1603 => x"94",
          1604 => x"cc",
          1605 => x"d9",
          1606 => x"80",
          1607 => x"82",
          1608 => x"43",
          1609 => x"84",
          1610 => x"78",
          1611 => x"38",
          1612 => x"08",
          1613 => x"82",
          1614 => x"59",
          1615 => x"88",
          1616 => x"ac",
          1617 => x"39",
          1618 => x"33",
          1619 => x"2e",
          1620 => x"84",
          1621 => x"88",
          1622 => x"c0",
          1623 => x"43",
          1624 => x"f8",
          1625 => x"84",
          1626 => x"e9",
          1627 => x"ec",
          1628 => x"a9",
          1629 => x"5c",
          1630 => x"2e",
          1631 => x"5c",
          1632 => x"70",
          1633 => x"70",
          1634 => x"2a",
          1635 => x"51",
          1636 => x"78",
          1637 => x"38",
          1638 => x"83",
          1639 => x"81",
          1640 => x"9b",
          1641 => x"55",
          1642 => x"53",
          1643 => x"51",
          1644 => x"81",
          1645 => x"9b",
          1646 => x"d8",
          1647 => x"ff",
          1648 => x"ff",
          1649 => x"a3",
          1650 => x"85",
          1651 => x"2e",
          1652 => x"b4",
          1653 => x"11",
          1654 => x"05",
          1655 => x"3f",
          1656 => x"08",
          1657 => x"38",
          1658 => x"80",
          1659 => x"79",
          1660 => x"05",
          1661 => x"fe",
          1662 => x"ff",
          1663 => x"a2",
          1664 => x"85",
          1665 => x"38",
          1666 => x"63",
          1667 => x"52",
          1668 => x"51",
          1669 => x"80",
          1670 => x"51",
          1671 => x"79",
          1672 => x"59",
          1673 => x"f8",
          1674 => x"79",
          1675 => x"b4",
          1676 => x"11",
          1677 => x"05",
          1678 => x"3f",
          1679 => x"08",
          1680 => x"38",
          1681 => x"80",
          1682 => x"79",
          1683 => x"05",
          1684 => x"39",
          1685 => x"51",
          1686 => x"ff",
          1687 => x"3d",
          1688 => x"53",
          1689 => x"51",
          1690 => x"82",
          1691 => x"80",
          1692 => x"38",
          1693 => x"f0",
          1694 => x"84",
          1695 => x"d1",
          1696 => x"ec",
          1697 => x"a5",
          1698 => x"02",
          1699 => x"79",
          1700 => x"5b",
          1701 => x"b4",
          1702 => x"11",
          1703 => x"05",
          1704 => x"3f",
          1705 => x"08",
          1706 => x"e8",
          1707 => x"22",
          1708 => x"f3",
          1709 => x"a5",
          1710 => x"52",
          1711 => x"f7",
          1712 => x"79",
          1713 => x"ae",
          1714 => x"38",
          1715 => x"87",
          1716 => x"05",
          1717 => x"b4",
          1718 => x"11",
          1719 => x"05",
          1720 => x"3f",
          1721 => x"08",
          1722 => x"38",
          1723 => x"be",
          1724 => x"70",
          1725 => x"23",
          1726 => x"b1",
          1727 => x"84",
          1728 => x"3f",
          1729 => x"b4",
          1730 => x"11",
          1731 => x"05",
          1732 => x"3f",
          1733 => x"08",
          1734 => x"f8",
          1735 => x"fe",
          1736 => x"ff",
          1737 => x"a2",
          1738 => x"85",
          1739 => x"2e",
          1740 => x"60",
          1741 => x"60",
          1742 => x"b4",
          1743 => x"11",
          1744 => x"05",
          1745 => x"3f",
          1746 => x"08",
          1747 => x"c4",
          1748 => x"08",
          1749 => x"f3",
          1750 => x"81",
          1751 => x"52",
          1752 => x"d3",
          1753 => x"79",
          1754 => x"ae",
          1755 => x"38",
          1756 => x"9b",
          1757 => x"fe",
          1758 => x"ff",
          1759 => x"a1",
          1760 => x"85",
          1761 => x"2e",
          1762 => x"60",
          1763 => x"60",
          1764 => x"ff",
          1765 => x"f3",
          1766 => x"d1",
          1767 => x"39",
          1768 => x"80",
          1769 => x"84",
          1770 => x"a9",
          1771 => x"ec",
          1772 => x"f5",
          1773 => x"52",
          1774 => x"51",
          1775 => x"63",
          1776 => x"b4",
          1777 => x"11",
          1778 => x"05",
          1779 => x"3f",
          1780 => x"08",
          1781 => x"bc",
          1782 => x"81",
          1783 => x"9c",
          1784 => x"59",
          1785 => x"85",
          1786 => x"2e",
          1787 => x"82",
          1788 => x"52",
          1789 => x"51",
          1790 => x"f5",
          1791 => x"f3",
          1792 => x"e9",
          1793 => x"3f",
          1794 => x"81",
          1795 => x"96",
          1796 => x"59",
          1797 => x"90",
          1798 => x"f8",
          1799 => x"79",
          1800 => x"80",
          1801 => x"38",
          1802 => x"59",
          1803 => x"81",
          1804 => x"3d",
          1805 => x"51",
          1806 => x"82",
          1807 => x"5c",
          1808 => x"82",
          1809 => x"7a",
          1810 => x"38",
          1811 => x"8c",
          1812 => x"39",
          1813 => x"ae",
          1814 => x"39",
          1815 => x"56",
          1816 => x"f4",
          1817 => x"53",
          1818 => x"52",
          1819 => x"b0",
          1820 => x"ff",
          1821 => x"81",
          1822 => x"b4",
          1823 => x"05",
          1824 => x"3f",
          1825 => x"55",
          1826 => x"54",
          1827 => x"f4",
          1828 => x"3d",
          1829 => x"51",
          1830 => x"92",
          1831 => x"80",
          1832 => x"cc",
          1833 => x"ff",
          1834 => x"9b",
          1835 => x"84",
          1836 => x"85",
          1837 => x"56",
          1838 => x"54",
          1839 => x"53",
          1840 => x"52",
          1841 => x"b0",
          1842 => x"dc",
          1843 => x"ec",
          1844 => x"ec",
          1845 => x"09",
          1846 => x"72",
          1847 => x"51",
          1848 => x"80",
          1849 => x"26",
          1850 => x"5a",
          1851 => x"59",
          1852 => x"8d",
          1853 => x"70",
          1854 => x"5c",
          1855 => x"c2",
          1856 => x"32",
          1857 => x"07",
          1858 => x"38",
          1859 => x"09",
          1860 => x"80",
          1861 => x"d4",
          1862 => x"3f",
          1863 => x"fc",
          1864 => x"0b",
          1865 => x"34",
          1866 => x"8c",
          1867 => x"55",
          1868 => x"52",
          1869 => x"d4",
          1870 => x"ec",
          1871 => x"75",
          1872 => x"87",
          1873 => x"73",
          1874 => x"3f",
          1875 => x"ec",
          1876 => x"0c",
          1877 => x"9c",
          1878 => x"55",
          1879 => x"52",
          1880 => x"a8",
          1881 => x"ec",
          1882 => x"75",
          1883 => x"87",
          1884 => x"73",
          1885 => x"3f",
          1886 => x"ec",
          1887 => x"0c",
          1888 => x"0b",
          1889 => x"84",
          1890 => x"83",
          1891 => x"94",
          1892 => x"c0",
          1893 => x"9c",
          1894 => x"c3",
          1895 => x"9c",
          1896 => x"98",
          1897 => x"3f",
          1898 => x"51",
          1899 => x"81",
          1900 => x"93",
          1901 => x"85",
          1902 => x"3f",
          1903 => x"8c",
          1904 => x"3f",
          1905 => x"3d",
          1906 => x"83",
          1907 => x"2b",
          1908 => x"3f",
          1909 => x"08",
          1910 => x"72",
          1911 => x"54",
          1912 => x"25",
          1913 => x"82",
          1914 => x"84",
          1915 => x"fc",
          1916 => x"70",
          1917 => x"80",
          1918 => x"72",
          1919 => x"8c",
          1920 => x"51",
          1921 => x"09",
          1922 => x"38",
          1923 => x"f1",
          1924 => x"51",
          1925 => x"09",
          1926 => x"38",
          1927 => x"81",
          1928 => x"73",
          1929 => x"81",
          1930 => x"84",
          1931 => x"52",
          1932 => x"52",
          1933 => x"2e",
          1934 => x"54",
          1935 => x"9d",
          1936 => x"38",
          1937 => x"12",
          1938 => x"33",
          1939 => x"a0",
          1940 => x"81",
          1941 => x"2e",
          1942 => x"ea",
          1943 => x"33",
          1944 => x"a0",
          1945 => x"06",
          1946 => x"54",
          1947 => x"70",
          1948 => x"70",
          1949 => x"07",
          1950 => x"70",
          1951 => x"38",
          1952 => x"81",
          1953 => x"71",
          1954 => x"51",
          1955 => x"ec",
          1956 => x"0d",
          1957 => x"0d",
          1958 => x"08",
          1959 => x"38",
          1960 => x"05",
          1961 => x"9b",
          1962 => x"85",
          1963 => x"38",
          1964 => x"39",
          1965 => x"82",
          1966 => x"86",
          1967 => x"fc",
          1968 => x"82",
          1969 => x"05",
          1970 => x"52",
          1971 => x"81",
          1972 => x"13",
          1973 => x"51",
          1974 => x"9e",
          1975 => x"38",
          1976 => x"51",
          1977 => x"97",
          1978 => x"38",
          1979 => x"51",
          1980 => x"bb",
          1981 => x"38",
          1982 => x"51",
          1983 => x"bb",
          1984 => x"38",
          1985 => x"55",
          1986 => x"87",
          1987 => x"d9",
          1988 => x"22",
          1989 => x"73",
          1990 => x"80",
          1991 => x"0b",
          1992 => x"9c",
          1993 => x"87",
          1994 => x"0c",
          1995 => x"87",
          1996 => x"0c",
          1997 => x"87",
          1998 => x"0c",
          1999 => x"87",
          2000 => x"0c",
          2001 => x"87",
          2002 => x"0c",
          2003 => x"87",
          2004 => x"0c",
          2005 => x"98",
          2006 => x"87",
          2007 => x"0c",
          2008 => x"c0",
          2009 => x"80",
          2010 => x"85",
          2011 => x"3d",
          2012 => x"3d",
          2013 => x"87",
          2014 => x"5d",
          2015 => x"87",
          2016 => x"08",
          2017 => x"23",
          2018 => x"b8",
          2019 => x"82",
          2020 => x"c0",
          2021 => x"5a",
          2022 => x"34",
          2023 => x"b0",
          2024 => x"84",
          2025 => x"c0",
          2026 => x"5a",
          2027 => x"34",
          2028 => x"a8",
          2029 => x"86",
          2030 => x"c0",
          2031 => x"5c",
          2032 => x"23",
          2033 => x"a0",
          2034 => x"8a",
          2035 => x"7d",
          2036 => x"ff",
          2037 => x"7b",
          2038 => x"06",
          2039 => x"33",
          2040 => x"33",
          2041 => x"33",
          2042 => x"33",
          2043 => x"33",
          2044 => x"ff",
          2045 => x"81",
          2046 => x"94",
          2047 => x"3d",
          2048 => x"3d",
          2049 => x"05",
          2050 => x"81",
          2051 => x"2a",
          2052 => x"70",
          2053 => x"34",
          2054 => x"04",
          2055 => x"77",
          2056 => x"33",
          2057 => x"06",
          2058 => x"87",
          2059 => x"51",
          2060 => x"86",
          2061 => x"94",
          2062 => x"08",
          2063 => x"70",
          2064 => x"54",
          2065 => x"2e",
          2066 => x"91",
          2067 => x"06",
          2068 => x"d7",
          2069 => x"32",
          2070 => x"51",
          2071 => x"2e",
          2072 => x"93",
          2073 => x"06",
          2074 => x"ff",
          2075 => x"81",
          2076 => x"87",
          2077 => x"52",
          2078 => x"86",
          2079 => x"94",
          2080 => x"72",
          2081 => x"85",
          2082 => x"3d",
          2083 => x"3d",
          2084 => x"05",
          2085 => x"8c",
          2086 => x"ff",
          2087 => x"56",
          2088 => x"84",
          2089 => x"2e",
          2090 => x"c0",
          2091 => x"70",
          2092 => x"2a",
          2093 => x"53",
          2094 => x"80",
          2095 => x"71",
          2096 => x"81",
          2097 => x"70",
          2098 => x"81",
          2099 => x"06",
          2100 => x"80",
          2101 => x"71",
          2102 => x"81",
          2103 => x"70",
          2104 => x"73",
          2105 => x"51",
          2106 => x"80",
          2107 => x"2e",
          2108 => x"c0",
          2109 => x"75",
          2110 => x"3d",
          2111 => x"3d",
          2112 => x"80",
          2113 => x"81",
          2114 => x"53",
          2115 => x"2e",
          2116 => x"71",
          2117 => x"81",
          2118 => x"8c",
          2119 => x"ff",
          2120 => x"55",
          2121 => x"94",
          2122 => x"80",
          2123 => x"87",
          2124 => x"51",
          2125 => x"96",
          2126 => x"06",
          2127 => x"70",
          2128 => x"38",
          2129 => x"70",
          2130 => x"51",
          2131 => x"72",
          2132 => x"81",
          2133 => x"70",
          2134 => x"38",
          2135 => x"70",
          2136 => x"51",
          2137 => x"38",
          2138 => x"06",
          2139 => x"94",
          2140 => x"80",
          2141 => x"87",
          2142 => x"52",
          2143 => x"81",
          2144 => x"70",
          2145 => x"53",
          2146 => x"ff",
          2147 => x"82",
          2148 => x"89",
          2149 => x"fe",
          2150 => x"84",
          2151 => x"81",
          2152 => x"52",
          2153 => x"84",
          2154 => x"2e",
          2155 => x"c0",
          2156 => x"70",
          2157 => x"2a",
          2158 => x"51",
          2159 => x"80",
          2160 => x"71",
          2161 => x"51",
          2162 => x"80",
          2163 => x"2e",
          2164 => x"c0",
          2165 => x"71",
          2166 => x"ff",
          2167 => x"ec",
          2168 => x"3d",
          2169 => x"3d",
          2170 => x"8c",
          2171 => x"ff",
          2172 => x"87",
          2173 => x"52",
          2174 => x"86",
          2175 => x"94",
          2176 => x"08",
          2177 => x"70",
          2178 => x"51",
          2179 => x"70",
          2180 => x"38",
          2181 => x"06",
          2182 => x"94",
          2183 => x"80",
          2184 => x"87",
          2185 => x"52",
          2186 => x"98",
          2187 => x"2c",
          2188 => x"71",
          2189 => x"0c",
          2190 => x"04",
          2191 => x"87",
          2192 => x"08",
          2193 => x"8a",
          2194 => x"70",
          2195 => x"b4",
          2196 => x"9e",
          2197 => x"84",
          2198 => x"c0",
          2199 => x"82",
          2200 => x"87",
          2201 => x"08",
          2202 => x"0c",
          2203 => x"98",
          2204 => x"9c",
          2205 => x"9e",
          2206 => x"84",
          2207 => x"c0",
          2208 => x"82",
          2209 => x"87",
          2210 => x"08",
          2211 => x"0c",
          2212 => x"b0",
          2213 => x"ac",
          2214 => x"9e",
          2215 => x"84",
          2216 => x"c0",
          2217 => x"82",
          2218 => x"87",
          2219 => x"08",
          2220 => x"0c",
          2221 => x"c0",
          2222 => x"bc",
          2223 => x"9e",
          2224 => x"84",
          2225 => x"c0",
          2226 => x"51",
          2227 => x"c4",
          2228 => x"9e",
          2229 => x"84",
          2230 => x"c0",
          2231 => x"82",
          2232 => x"87",
          2233 => x"08",
          2234 => x"0c",
          2235 => x"84",
          2236 => x"0b",
          2237 => x"90",
          2238 => x"80",
          2239 => x"52",
          2240 => x"2e",
          2241 => x"52",
          2242 => x"d5",
          2243 => x"87",
          2244 => x"08",
          2245 => x"0a",
          2246 => x"52",
          2247 => x"83",
          2248 => x"71",
          2249 => x"34",
          2250 => x"c0",
          2251 => x"70",
          2252 => x"06",
          2253 => x"70",
          2254 => x"38",
          2255 => x"82",
          2256 => x"80",
          2257 => x"9e",
          2258 => x"88",
          2259 => x"51",
          2260 => x"80",
          2261 => x"81",
          2262 => x"84",
          2263 => x"0b",
          2264 => x"90",
          2265 => x"80",
          2266 => x"52",
          2267 => x"2e",
          2268 => x"52",
          2269 => x"d9",
          2270 => x"87",
          2271 => x"08",
          2272 => x"80",
          2273 => x"52",
          2274 => x"83",
          2275 => x"71",
          2276 => x"34",
          2277 => x"c0",
          2278 => x"70",
          2279 => x"06",
          2280 => x"70",
          2281 => x"38",
          2282 => x"82",
          2283 => x"80",
          2284 => x"9e",
          2285 => x"82",
          2286 => x"51",
          2287 => x"80",
          2288 => x"81",
          2289 => x"84",
          2290 => x"0b",
          2291 => x"90",
          2292 => x"80",
          2293 => x"52",
          2294 => x"2e",
          2295 => x"52",
          2296 => x"dd",
          2297 => x"87",
          2298 => x"08",
          2299 => x"80",
          2300 => x"52",
          2301 => x"83",
          2302 => x"71",
          2303 => x"34",
          2304 => x"c0",
          2305 => x"70",
          2306 => x"51",
          2307 => x"80",
          2308 => x"81",
          2309 => x"84",
          2310 => x"c0",
          2311 => x"70",
          2312 => x"70",
          2313 => x"51",
          2314 => x"84",
          2315 => x"0b",
          2316 => x"90",
          2317 => x"80",
          2318 => x"52",
          2319 => x"83",
          2320 => x"71",
          2321 => x"34",
          2322 => x"90",
          2323 => x"f0",
          2324 => x"2a",
          2325 => x"70",
          2326 => x"34",
          2327 => x"c0",
          2328 => x"70",
          2329 => x"52",
          2330 => x"2e",
          2331 => x"52",
          2332 => x"e3",
          2333 => x"9e",
          2334 => x"87",
          2335 => x"70",
          2336 => x"34",
          2337 => x"04",
          2338 => x"81",
          2339 => x"85",
          2340 => x"84",
          2341 => x"73",
          2342 => x"38",
          2343 => x"51",
          2344 => x"81",
          2345 => x"85",
          2346 => x"84",
          2347 => x"73",
          2348 => x"38",
          2349 => x"08",
          2350 => x"08",
          2351 => x"81",
          2352 => x"8b",
          2353 => x"84",
          2354 => x"73",
          2355 => x"38",
          2356 => x"08",
          2357 => x"08",
          2358 => x"81",
          2359 => x"8a",
          2360 => x"84",
          2361 => x"73",
          2362 => x"38",
          2363 => x"08",
          2364 => x"08",
          2365 => x"81",
          2366 => x"8a",
          2367 => x"84",
          2368 => x"73",
          2369 => x"38",
          2370 => x"08",
          2371 => x"08",
          2372 => x"81",
          2373 => x"8a",
          2374 => x"84",
          2375 => x"73",
          2376 => x"38",
          2377 => x"08",
          2378 => x"08",
          2379 => x"81",
          2380 => x"8a",
          2381 => x"84",
          2382 => x"73",
          2383 => x"38",
          2384 => x"33",
          2385 => x"ec",
          2386 => x"3f",
          2387 => x"33",
          2388 => x"2e",
          2389 => x"84",
          2390 => x"81",
          2391 => x"89",
          2392 => x"84",
          2393 => x"73",
          2394 => x"38",
          2395 => x"33",
          2396 => x"ac",
          2397 => x"3f",
          2398 => x"33",
          2399 => x"2e",
          2400 => x"f7",
          2401 => x"e5",
          2402 => x"d7",
          2403 => x"80",
          2404 => x"81",
          2405 => x"83",
          2406 => x"84",
          2407 => x"73",
          2408 => x"38",
          2409 => x"51",
          2410 => x"82",
          2411 => x"54",
          2412 => x"88",
          2413 => x"f8",
          2414 => x"3f",
          2415 => x"33",
          2416 => x"2e",
          2417 => x"f8",
          2418 => x"a1",
          2419 => x"90",
          2420 => x"3f",
          2421 => x"08",
          2422 => x"9c",
          2423 => x"3f",
          2424 => x"08",
          2425 => x"c4",
          2426 => x"3f",
          2427 => x"08",
          2428 => x"ec",
          2429 => x"3f",
          2430 => x"51",
          2431 => x"82",
          2432 => x"52",
          2433 => x"51",
          2434 => x"82",
          2435 => x"55",
          2436 => x"52",
          2437 => x"f4",
          2438 => x"ec",
          2439 => x"84",
          2440 => x"85",
          2441 => x"d0",
          2442 => x"82",
          2443 => x"31",
          2444 => x"81",
          2445 => x"88",
          2446 => x"84",
          2447 => x"73",
          2448 => x"38",
          2449 => x"08",
          2450 => x"c0",
          2451 => x"d1",
          2452 => x"85",
          2453 => x"bd",
          2454 => x"82",
          2455 => x"51",
          2456 => x"74",
          2457 => x"08",
          2458 => x"52",
          2459 => x"51",
          2460 => x"82",
          2461 => x"54",
          2462 => x"b0",
          2463 => x"d0",
          2464 => x"84",
          2465 => x"51",
          2466 => x"82",
          2467 => x"54",
          2468 => x"52",
          2469 => x"08",
          2470 => x"3f",
          2471 => x"ec",
          2472 => x"73",
          2473 => x"9c",
          2474 => x"3f",
          2475 => x"51",
          2476 => x"86",
          2477 => x"fe",
          2478 => x"92",
          2479 => x"05",
          2480 => x"26",
          2481 => x"82",
          2482 => x"e8",
          2483 => x"04",
          2484 => x"51",
          2485 => x"fa",
          2486 => x"39",
          2487 => x"51",
          2488 => x"fa",
          2489 => x"39",
          2490 => x"51",
          2491 => x"fa",
          2492 => x"f9",
          2493 => x"0d",
          2494 => x"80",
          2495 => x"0b",
          2496 => x"84",
          2497 => x"84",
          2498 => x"c0",
          2499 => x"04",
          2500 => x"02",
          2501 => x"53",
          2502 => x"09",
          2503 => x"38",
          2504 => x"3f",
          2505 => x"08",
          2506 => x"2e",
          2507 => x"72",
          2508 => x"fc",
          2509 => x"82",
          2510 => x"8f",
          2511 => x"f4",
          2512 => x"80",
          2513 => x"72",
          2514 => x"84",
          2515 => x"fe",
          2516 => x"97",
          2517 => x"9c",
          2518 => x"82",
          2519 => x"54",
          2520 => x"3f",
          2521 => x"f4",
          2522 => x"0d",
          2523 => x"0d",
          2524 => x"33",
          2525 => x"06",
          2526 => x"80",
          2527 => x"72",
          2528 => x"51",
          2529 => x"ff",
          2530 => x"39",
          2531 => x"04",
          2532 => x"77",
          2533 => x"08",
          2534 => x"f4",
          2535 => x"73",
          2536 => x"ff",
          2537 => x"71",
          2538 => x"38",
          2539 => x"06",
          2540 => x"54",
          2541 => x"e7",
          2542 => x"9c",
          2543 => x"3d",
          2544 => x"3d",
          2545 => x"59",
          2546 => x"81",
          2547 => x"56",
          2548 => x"85",
          2549 => x"a5",
          2550 => x"06",
          2551 => x"80",
          2552 => x"81",
          2553 => x"58",
          2554 => x"b0",
          2555 => x"06",
          2556 => x"5a",
          2557 => x"ad",
          2558 => x"06",
          2559 => x"5a",
          2560 => x"05",
          2561 => x"75",
          2562 => x"81",
          2563 => x"77",
          2564 => x"08",
          2565 => x"05",
          2566 => x"5d",
          2567 => x"39",
          2568 => x"72",
          2569 => x"38",
          2570 => x"7b",
          2571 => x"18",
          2572 => x"70",
          2573 => x"33",
          2574 => x"53",
          2575 => x"80",
          2576 => x"09",
          2577 => x"72",
          2578 => x"78",
          2579 => x"70",
          2580 => x"70",
          2581 => x"25",
          2582 => x"54",
          2583 => x"53",
          2584 => x"8c",
          2585 => x"07",
          2586 => x"05",
          2587 => x"5a",
          2588 => x"83",
          2589 => x"54",
          2590 => x"27",
          2591 => x"16",
          2592 => x"06",
          2593 => x"80",
          2594 => x"aa",
          2595 => x"cf",
          2596 => x"73",
          2597 => x"81",
          2598 => x"80",
          2599 => x"38",
          2600 => x"2e",
          2601 => x"81",
          2602 => x"80",
          2603 => x"8a",
          2604 => x"39",
          2605 => x"2e",
          2606 => x"73",
          2607 => x"8a",
          2608 => x"d3",
          2609 => x"80",
          2610 => x"80",
          2611 => x"ee",
          2612 => x"39",
          2613 => x"71",
          2614 => x"53",
          2615 => x"54",
          2616 => x"2e",
          2617 => x"15",
          2618 => x"33",
          2619 => x"72",
          2620 => x"81",
          2621 => x"39",
          2622 => x"56",
          2623 => x"27",
          2624 => x"51",
          2625 => x"75",
          2626 => x"72",
          2627 => x"38",
          2628 => x"d9",
          2629 => x"16",
          2630 => x"7b",
          2631 => x"38",
          2632 => x"ec",
          2633 => x"77",
          2634 => x"12",
          2635 => x"53",
          2636 => x"5c",
          2637 => x"5c",
          2638 => x"5c",
          2639 => x"5c",
          2640 => x"51",
          2641 => x"fd",
          2642 => x"82",
          2643 => x"06",
          2644 => x"80",
          2645 => x"77",
          2646 => x"53",
          2647 => x"18",
          2648 => x"72",
          2649 => x"c4",
          2650 => x"81",
          2651 => x"07",
          2652 => x"55",
          2653 => x"80",
          2654 => x"72",
          2655 => x"38",
          2656 => x"05",
          2657 => x"5b",
          2658 => x"8f",
          2659 => x"7b",
          2660 => x"cb",
          2661 => x"85",
          2662 => x"ff",
          2663 => x"75",
          2664 => x"e8",
          2665 => x"ec",
          2666 => x"74",
          2667 => x"a7",
          2668 => x"80",
          2669 => x"38",
          2670 => x"72",
          2671 => x"54",
          2672 => x"72",
          2673 => x"05",
          2674 => x"17",
          2675 => x"05",
          2676 => x"9f",
          2677 => x"57",
          2678 => x"85",
          2679 => x"af",
          2680 => x"2a",
          2681 => x"51",
          2682 => x"2e",
          2683 => x"3d",
          2684 => x"05",
          2685 => x"34",
          2686 => x"76",
          2687 => x"54",
          2688 => x"72",
          2689 => x"54",
          2690 => x"70",
          2691 => x"56",
          2692 => x"81",
          2693 => x"7b",
          2694 => x"73",
          2695 => x"3f",
          2696 => x"53",
          2697 => x"74",
          2698 => x"53",
          2699 => x"eb",
          2700 => x"77",
          2701 => x"53",
          2702 => x"14",
          2703 => x"54",
          2704 => x"3f",
          2705 => x"74",
          2706 => x"53",
          2707 => x"fa",
          2708 => x"51",
          2709 => x"ef",
          2710 => x"0d",
          2711 => x"0d",
          2712 => x"70",
          2713 => x"08",
          2714 => x"51",
          2715 => x"85",
          2716 => x"fe",
          2717 => x"82",
          2718 => x"85",
          2719 => x"52",
          2720 => x"be",
          2721 => x"fc",
          2722 => x"73",
          2723 => x"82",
          2724 => x"84",
          2725 => x"fd",
          2726 => x"9c",
          2727 => x"82",
          2728 => x"87",
          2729 => x"53",
          2730 => x"fa",
          2731 => x"82",
          2732 => x"85",
          2733 => x"fb",
          2734 => x"79",
          2735 => x"08",
          2736 => x"57",
          2737 => x"71",
          2738 => x"e3",
          2739 => x"f8",
          2740 => x"2d",
          2741 => x"08",
          2742 => x"53",
          2743 => x"80",
          2744 => x"8d",
          2745 => x"72",
          2746 => x"09",
          2747 => x"80",
          2748 => x"52",
          2749 => x"8b",
          2750 => x"2e",
          2751 => x"14",
          2752 => x"9f",
          2753 => x"38",
          2754 => x"73",
          2755 => x"bd",
          2756 => x"52",
          2757 => x"81",
          2758 => x"51",
          2759 => x"ff",
          2760 => x"15",
          2761 => x"34",
          2762 => x"e4",
          2763 => x"72",
          2764 => x"0c",
          2765 => x"04",
          2766 => x"82",
          2767 => x"75",
          2768 => x"0c",
          2769 => x"52",
          2770 => x"3f",
          2771 => x"f8",
          2772 => x"0d",
          2773 => x"0d",
          2774 => x"56",
          2775 => x"0c",
          2776 => x"70",
          2777 => x"73",
          2778 => x"81",
          2779 => x"81",
          2780 => x"ed",
          2781 => x"2e",
          2782 => x"8e",
          2783 => x"08",
          2784 => x"76",
          2785 => x"56",
          2786 => x"b0",
          2787 => x"06",
          2788 => x"75",
          2789 => x"76",
          2790 => x"70",
          2791 => x"73",
          2792 => x"8b",
          2793 => x"73",
          2794 => x"85",
          2795 => x"82",
          2796 => x"76",
          2797 => x"70",
          2798 => x"ac",
          2799 => x"a0",
          2800 => x"84",
          2801 => x"53",
          2802 => x"57",
          2803 => x"98",
          2804 => x"39",
          2805 => x"80",
          2806 => x"26",
          2807 => x"86",
          2808 => x"80",
          2809 => x"57",
          2810 => x"74",
          2811 => x"38",
          2812 => x"27",
          2813 => x"14",
          2814 => x"06",
          2815 => x"14",
          2816 => x"06",
          2817 => x"74",
          2818 => x"f9",
          2819 => x"ff",
          2820 => x"89",
          2821 => x"38",
          2822 => x"c5",
          2823 => x"74",
          2824 => x"3f",
          2825 => x"08",
          2826 => x"81",
          2827 => x"76",
          2828 => x"56",
          2829 => x"b2",
          2830 => x"2e",
          2831 => x"09",
          2832 => x"74",
          2833 => x"55",
          2834 => x"ec",
          2835 => x"0d",
          2836 => x"0d",
          2837 => x"56",
          2838 => x"0c",
          2839 => x"70",
          2840 => x"73",
          2841 => x"81",
          2842 => x"81",
          2843 => x"ed",
          2844 => x"2e",
          2845 => x"8e",
          2846 => x"08",
          2847 => x"76",
          2848 => x"56",
          2849 => x"b0",
          2850 => x"06",
          2851 => x"75",
          2852 => x"76",
          2853 => x"70",
          2854 => x"73",
          2855 => x"8b",
          2856 => x"73",
          2857 => x"85",
          2858 => x"82",
          2859 => x"76",
          2860 => x"70",
          2861 => x"ac",
          2862 => x"a0",
          2863 => x"84",
          2864 => x"53",
          2865 => x"57",
          2866 => x"98",
          2867 => x"39",
          2868 => x"80",
          2869 => x"26",
          2870 => x"86",
          2871 => x"80",
          2872 => x"57",
          2873 => x"74",
          2874 => x"38",
          2875 => x"27",
          2876 => x"14",
          2877 => x"06",
          2878 => x"14",
          2879 => x"06",
          2880 => x"74",
          2881 => x"f9",
          2882 => x"ff",
          2883 => x"89",
          2884 => x"38",
          2885 => x"c5",
          2886 => x"74",
          2887 => x"3f",
          2888 => x"08",
          2889 => x"81",
          2890 => x"76",
          2891 => x"56",
          2892 => x"b2",
          2893 => x"2e",
          2894 => x"09",
          2895 => x"74",
          2896 => x"55",
          2897 => x"ec",
          2898 => x"0d",
          2899 => x"0d",
          2900 => x"70",
          2901 => x"98",
          2902 => x"2c",
          2903 => x"11",
          2904 => x"56",
          2905 => x"51",
          2906 => x"fa",
          2907 => x"55",
          2908 => x"25",
          2909 => x"81",
          2910 => x"08",
          2911 => x"05",
          2912 => x"71",
          2913 => x"53",
          2914 => x"2e",
          2915 => x"83",
          2916 => x"73",
          2917 => x"85",
          2918 => x"3d",
          2919 => x"3d",
          2920 => x"84",
          2921 => x"33",
          2922 => x"55",
          2923 => x"2e",
          2924 => x"51",
          2925 => x"a0",
          2926 => x"3f",
          2927 => x"d0",
          2928 => x"ff",
          2929 => x"73",
          2930 => x"ff",
          2931 => x"39",
          2932 => x"99",
          2933 => x"34",
          2934 => x"04",
          2935 => x"7c",
          2936 => x"b7",
          2937 => x"88",
          2938 => x"33",
          2939 => x"33",
          2940 => x"82",
          2941 => x"08",
          2942 => x"5a",
          2943 => x"80",
          2944 => x"74",
          2945 => x"3f",
          2946 => x"33",
          2947 => x"82",
          2948 => x"81",
          2949 => x"59",
          2950 => x"9d",
          2951 => x"85",
          2952 => x"0c",
          2953 => x"33",
          2954 => x"82",
          2955 => x"08",
          2956 => x"74",
          2957 => x"38",
          2958 => x"52",
          2959 => x"b8",
          2960 => x"85",
          2961 => x"05",
          2962 => x"85",
          2963 => x"81",
          2964 => x"93",
          2965 => x"38",
          2966 => x"85",
          2967 => x"80",
          2968 => x"82",
          2969 => x"56",
          2970 => x"ac",
          2971 => x"bc",
          2972 => x"a4",
          2973 => x"fc",
          2974 => x"53",
          2975 => x"51",
          2976 => x"3f",
          2977 => x"08",
          2978 => x"81",
          2979 => x"82",
          2980 => x"51",
          2981 => x"3f",
          2982 => x"04",
          2983 => x"82",
          2984 => x"93",
          2985 => x"52",
          2986 => x"89",
          2987 => x"98",
          2988 => x"73",
          2989 => x"84",
          2990 => x"73",
          2991 => x"38",
          2992 => x"85",
          2993 => x"85",
          2994 => x"71",
          2995 => x"38",
          2996 => x"d9",
          2997 => x"85",
          2998 => x"98",
          2999 => x"0b",
          3000 => x"0c",
          3001 => x"04",
          3002 => x"81",
          3003 => x"82",
          3004 => x"51",
          3005 => x"3f",
          3006 => x"08",
          3007 => x"82",
          3008 => x"53",
          3009 => x"88",
          3010 => x"56",
          3011 => x"3f",
          3012 => x"08",
          3013 => x"38",
          3014 => x"b5",
          3015 => x"85",
          3016 => x"80",
          3017 => x"ec",
          3018 => x"38",
          3019 => x"08",
          3020 => x"17",
          3021 => x"74",
          3022 => x"76",
          3023 => x"81",
          3024 => x"57",
          3025 => x"74",
          3026 => x"81",
          3027 => x"38",
          3028 => x"04",
          3029 => x"aa",
          3030 => x"3d",
          3031 => x"81",
          3032 => x"80",
          3033 => x"c0",
          3034 => x"dd",
          3035 => x"85",
          3036 => x"96",
          3037 => x"82",
          3038 => x"54",
          3039 => x"52",
          3040 => x"52",
          3041 => x"ba",
          3042 => x"ec",
          3043 => x"a5",
          3044 => x"ff",
          3045 => x"82",
          3046 => x"81",
          3047 => x"80",
          3048 => x"ec",
          3049 => x"38",
          3050 => x"08",
          3051 => x"17",
          3052 => x"74",
          3053 => x"70",
          3054 => x"70",
          3055 => x"2a",
          3056 => x"78",
          3057 => x"38",
          3058 => x"38",
          3059 => x"08",
          3060 => x"53",
          3061 => x"e7",
          3062 => x"ec",
          3063 => x"88",
          3064 => x"f4",
          3065 => x"3f",
          3066 => x"09",
          3067 => x"38",
          3068 => x"51",
          3069 => x"3f",
          3070 => x"b3",
          3071 => x"3d",
          3072 => x"85",
          3073 => x"34",
          3074 => x"82",
          3075 => x"a9",
          3076 => x"f6",
          3077 => x"7e",
          3078 => x"72",
          3079 => x"5a",
          3080 => x"2e",
          3081 => x"a2",
          3082 => x"78",
          3083 => x"76",
          3084 => x"81",
          3085 => x"70",
          3086 => x"58",
          3087 => x"2e",
          3088 => x"86",
          3089 => x"26",
          3090 => x"55",
          3091 => x"82",
          3092 => x"70",
          3093 => x"54",
          3094 => x"3f",
          3095 => x"08",
          3096 => x"73",
          3097 => x"b5",
          3098 => x"85",
          3099 => x"c3",
          3100 => x"33",
          3101 => x"2e",
          3102 => x"82",
          3103 => x"b3",
          3104 => x"3f",
          3105 => x"1a",
          3106 => x"fc",
          3107 => x"05",
          3108 => x"3f",
          3109 => x"08",
          3110 => x"38",
          3111 => x"78",
          3112 => x"fd",
          3113 => x"85",
          3114 => x"ff",
          3115 => x"80",
          3116 => x"81",
          3117 => x"ff",
          3118 => x"82",
          3119 => x"8c",
          3120 => x"73",
          3121 => x"0c",
          3122 => x"04",
          3123 => x"b0",
          3124 => x"3d",
          3125 => x"08",
          3126 => x"80",
          3127 => x"34",
          3128 => x"33",
          3129 => x"08",
          3130 => x"81",
          3131 => x"82",
          3132 => x"55",
          3133 => x"38",
          3134 => x"80",
          3135 => x"38",
          3136 => x"06",
          3137 => x"80",
          3138 => x"38",
          3139 => x"95",
          3140 => x"ec",
          3141 => x"c0",
          3142 => x"ec",
          3143 => x"81",
          3144 => x"53",
          3145 => x"85",
          3146 => x"80",
          3147 => x"82",
          3148 => x"80",
          3149 => x"81",
          3150 => x"f2",
          3151 => x"f7",
          3152 => x"ec",
          3153 => x"85",
          3154 => x"80",
          3155 => x"3d",
          3156 => x"81",
          3157 => x"82",
          3158 => x"56",
          3159 => x"08",
          3160 => x"81",
          3161 => x"38",
          3162 => x"08",
          3163 => x"cb",
          3164 => x"ec",
          3165 => x"0b",
          3166 => x"08",
          3167 => x"82",
          3168 => x"ff",
          3169 => x"55",
          3170 => x"34",
          3171 => x"81",
          3172 => x"75",
          3173 => x"3f",
          3174 => x"81",
          3175 => x"54",
          3176 => x"83",
          3177 => x"74",
          3178 => x"81",
          3179 => x"38",
          3180 => x"82",
          3181 => x"76",
          3182 => x"85",
          3183 => x"2e",
          3184 => x"d8",
          3185 => x"5d",
          3186 => x"82",
          3187 => x"98",
          3188 => x"2c",
          3189 => x"ff",
          3190 => x"78",
          3191 => x"82",
          3192 => x"70",
          3193 => x"98",
          3194 => x"80",
          3195 => x"2b",
          3196 => x"71",
          3197 => x"70",
          3198 => x"fa",
          3199 => x"15",
          3200 => x"51",
          3201 => x"59",
          3202 => x"58",
          3203 => x"78",
          3204 => x"38",
          3205 => x"b1",
          3206 => x"70",
          3207 => x"98",
          3208 => x"54",
          3209 => x"80",
          3210 => x"53",
          3211 => x"51",
          3212 => x"82",
          3213 => x"81",
          3214 => x"73",
          3215 => x"38",
          3216 => x"80",
          3217 => x"ae",
          3218 => x"70",
          3219 => x"98",
          3220 => x"ff",
          3221 => x"56",
          3222 => x"26",
          3223 => x"53",
          3224 => x"51",
          3225 => x"82",
          3226 => x"81",
          3227 => x"73",
          3228 => x"39",
          3229 => x"80",
          3230 => x"38",
          3231 => x"73",
          3232 => x"34",
          3233 => x"70",
          3234 => x"9d",
          3235 => x"98",
          3236 => x"2c",
          3237 => x"11",
          3238 => x"fa",
          3239 => x"5e",
          3240 => x"58",
          3241 => x"73",
          3242 => x"81",
          3243 => x"38",
          3244 => x"15",
          3245 => x"80",
          3246 => x"84",
          3247 => x"82",
          3248 => x"92",
          3249 => x"9d",
          3250 => x"82",
          3251 => x"78",
          3252 => x"75",
          3253 => x"54",
          3254 => x"fd",
          3255 => x"82",
          3256 => x"e8",
          3257 => x"04",
          3258 => x"33",
          3259 => x"2e",
          3260 => x"82",
          3261 => x"54",
          3262 => x"ab",
          3263 => x"2b",
          3264 => x"51",
          3265 => x"24",
          3266 => x"1a",
          3267 => x"81",
          3268 => x"15",
          3269 => x"70",
          3270 => x"9d",
          3271 => x"51",
          3272 => x"74",
          3273 => x"82",
          3274 => x"81",
          3275 => x"74",
          3276 => x"34",
          3277 => x"ae",
          3278 => x"34",
          3279 => x"33",
          3280 => x"25",
          3281 => x"14",
          3282 => x"9d",
          3283 => x"9d",
          3284 => x"05",
          3285 => x"70",
          3286 => x"9d",
          3287 => x"51",
          3288 => x"76",
          3289 => x"74",
          3290 => x"52",
          3291 => x"3f",
          3292 => x"98",
          3293 => x"2c",
          3294 => x"33",
          3295 => x"54",
          3296 => x"e3",
          3297 => x"8c",
          3298 => x"2b",
          3299 => x"82",
          3300 => x"59",
          3301 => x"74",
          3302 => x"a9",
          3303 => x"e6",
          3304 => x"15",
          3305 => x"70",
          3306 => x"9d",
          3307 => x"51",
          3308 => x"75",
          3309 => x"fc",
          3310 => x"7a",
          3311 => x"81",
          3312 => x"9d",
          3313 => x"52",
          3314 => x"51",
          3315 => x"81",
          3316 => x"9d",
          3317 => x"81",
          3318 => x"55",
          3319 => x"fb",
          3320 => x"9d",
          3321 => x"05",
          3322 => x"9d",
          3323 => x"15",
          3324 => x"9d",
          3325 => x"51",
          3326 => x"82",
          3327 => x"70",
          3328 => x"98",
          3329 => x"88",
          3330 => x"56",
          3331 => x"25",
          3332 => x"1a",
          3333 => x"33",
          3334 => x"33",
          3335 => x"3f",
          3336 => x"98",
          3337 => x"2c",
          3338 => x"33",
          3339 => x"54",
          3340 => x"de",
          3341 => x"e5",
          3342 => x"9d",
          3343 => x"98",
          3344 => x"2c",
          3345 => x"33",
          3346 => x"57",
          3347 => x"fa",
          3348 => x"51",
          3349 => x"81",
          3350 => x"2b",
          3351 => x"82",
          3352 => x"59",
          3353 => x"75",
          3354 => x"38",
          3355 => x"82",
          3356 => x"7a",
          3357 => x"74",
          3358 => x"e5",
          3359 => x"9d",
          3360 => x"51",
          3361 => x"82",
          3362 => x"81",
          3363 => x"73",
          3364 => x"9d",
          3365 => x"73",
          3366 => x"38",
          3367 => x"52",
          3368 => x"b8",
          3369 => x"80",
          3370 => x"0b",
          3371 => x"34",
          3372 => x"9d",
          3373 => x"82",
          3374 => x"af",
          3375 => x"82",
          3376 => x"54",
          3377 => x"f9",
          3378 => x"51",
          3379 => x"82",
          3380 => x"ff",
          3381 => x"82",
          3382 => x"73",
          3383 => x"54",
          3384 => x"9d",
          3385 => x"9d",
          3386 => x"55",
          3387 => x"f9",
          3388 => x"14",
          3389 => x"9d",
          3390 => x"98",
          3391 => x"2c",
          3392 => x"06",
          3393 => x"74",
          3394 => x"38",
          3395 => x"81",
          3396 => x"34",
          3397 => x"e3",
          3398 => x"15",
          3399 => x"70",
          3400 => x"9d",
          3401 => x"51",
          3402 => x"75",
          3403 => x"a0",
          3404 => x"3f",
          3405 => x"33",
          3406 => x"70",
          3407 => x"9d",
          3408 => x"51",
          3409 => x"74",
          3410 => x"38",
          3411 => x"c0",
          3412 => x"70",
          3413 => x"98",
          3414 => x"88",
          3415 => x"56",
          3416 => x"25",
          3417 => x"dd",
          3418 => x"8c",
          3419 => x"ff",
          3420 => x"88",
          3421 => x"54",
          3422 => x"f8",
          3423 => x"14",
          3424 => x"9d",
          3425 => x"1a",
          3426 => x"54",
          3427 => x"82",
          3428 => x"70",
          3429 => x"82",
          3430 => x"58",
          3431 => x"75",
          3432 => x"f8",
          3433 => x"9d",
          3434 => x"52",
          3435 => x"51",
          3436 => x"80",
          3437 => x"8c",
          3438 => x"82",
          3439 => x"f8",
          3440 => x"b0",
          3441 => x"b8",
          3442 => x"80",
          3443 => x"74",
          3444 => x"e7",
          3445 => x"ec",
          3446 => x"88",
          3447 => x"ec",
          3448 => x"06",
          3449 => x"74",
          3450 => x"ff",
          3451 => x"93",
          3452 => x"39",
          3453 => x"82",
          3454 => x"fc",
          3455 => x"51",
          3456 => x"2e",
          3457 => x"51",
          3458 => x"3f",
          3459 => x"08",
          3460 => x"34",
          3461 => x"08",
          3462 => x"81",
          3463 => x"52",
          3464 => x"a8",
          3465 => x"1b",
          3466 => x"39",
          3467 => x"74",
          3468 => x"91",
          3469 => x"ff",
          3470 => x"99",
          3471 => x"2e",
          3472 => x"ae",
          3473 => x"ec",
          3474 => x"80",
          3475 => x"74",
          3476 => x"e7",
          3477 => x"ec",
          3478 => x"88",
          3479 => x"ec",
          3480 => x"06",
          3481 => x"74",
          3482 => x"ff",
          3483 => x"80",
          3484 => x"82",
          3485 => x"f0",
          3486 => x"54",
          3487 => x"ab",
          3488 => x"ff",
          3489 => x"82",
          3490 => x"82",
          3491 => x"82",
          3492 => x"81",
          3493 => x"05",
          3494 => x"79",
          3495 => x"fb",
          3496 => x"54",
          3497 => x"06",
          3498 => x"74",
          3499 => x"34",
          3500 => x"82",
          3501 => x"82",
          3502 => x"52",
          3503 => x"de",
          3504 => x"39",
          3505 => x"33",
          3506 => x"06",
          3507 => x"33",
          3508 => x"74",
          3509 => x"ed",
          3510 => x"54",
          3511 => x"8c",
          3512 => x"70",
          3513 => x"e0",
          3514 => x"d9",
          3515 => x"8c",
          3516 => x"80",
          3517 => x"38",
          3518 => x"94",
          3519 => x"8c",
          3520 => x"54",
          3521 => x"8c",
          3522 => x"39",
          3523 => x"83",
          3524 => x"82",
          3525 => x"82",
          3526 => x"85",
          3527 => x"80",
          3528 => x"83",
          3529 => x"ff",
          3530 => x"82",
          3531 => x"54",
          3532 => x"74",
          3533 => x"76",
          3534 => x"82",
          3535 => x"54",
          3536 => x"34",
          3537 => x"34",
          3538 => x"08",
          3539 => x"15",
          3540 => x"15",
          3541 => x"e4",
          3542 => x"e0",
          3543 => x"fe",
          3544 => x"70",
          3545 => x"06",
          3546 => x"58",
          3547 => x"74",
          3548 => x"73",
          3549 => x"82",
          3550 => x"70",
          3551 => x"85",
          3552 => x"f8",
          3553 => x"55",
          3554 => x"34",
          3555 => x"34",
          3556 => x"04",
          3557 => x"73",
          3558 => x"84",
          3559 => x"38",
          3560 => x"2a",
          3561 => x"83",
          3562 => x"51",
          3563 => x"82",
          3564 => x"83",
          3565 => x"f9",
          3566 => x"a6",
          3567 => x"84",
          3568 => x"22",
          3569 => x"85",
          3570 => x"83",
          3571 => x"74",
          3572 => x"11",
          3573 => x"12",
          3574 => x"2b",
          3575 => x"05",
          3576 => x"71",
          3577 => x"06",
          3578 => x"2a",
          3579 => x"59",
          3580 => x"57",
          3581 => x"71",
          3582 => x"81",
          3583 => x"85",
          3584 => x"75",
          3585 => x"54",
          3586 => x"34",
          3587 => x"34",
          3588 => x"08",
          3589 => x"33",
          3590 => x"71",
          3591 => x"70",
          3592 => x"ff",
          3593 => x"52",
          3594 => x"05",
          3595 => x"ff",
          3596 => x"2a",
          3597 => x"71",
          3598 => x"72",
          3599 => x"53",
          3600 => x"34",
          3601 => x"08",
          3602 => x"76",
          3603 => x"17",
          3604 => x"0d",
          3605 => x"0d",
          3606 => x"08",
          3607 => x"9e",
          3608 => x"83",
          3609 => x"86",
          3610 => x"12",
          3611 => x"2b",
          3612 => x"07",
          3613 => x"52",
          3614 => x"05",
          3615 => x"85",
          3616 => x"88",
          3617 => x"88",
          3618 => x"56",
          3619 => x"13",
          3620 => x"13",
          3621 => x"e4",
          3622 => x"84",
          3623 => x"12",
          3624 => x"2b",
          3625 => x"07",
          3626 => x"52",
          3627 => x"12",
          3628 => x"33",
          3629 => x"07",
          3630 => x"54",
          3631 => x"70",
          3632 => x"73",
          3633 => x"82",
          3634 => x"13",
          3635 => x"12",
          3636 => x"2b",
          3637 => x"ff",
          3638 => x"88",
          3639 => x"53",
          3640 => x"73",
          3641 => x"14",
          3642 => x"0d",
          3643 => x"0d",
          3644 => x"22",
          3645 => x"08",
          3646 => x"71",
          3647 => x"81",
          3648 => x"88",
          3649 => x"83",
          3650 => x"5b",
          3651 => x"05",
          3652 => x"12",
          3653 => x"2b",
          3654 => x"07",
          3655 => x"53",
          3656 => x"25",
          3657 => x"73",
          3658 => x"3f",
          3659 => x"08",
          3660 => x"33",
          3661 => x"71",
          3662 => x"83",
          3663 => x"11",
          3664 => x"12",
          3665 => x"2b",
          3666 => x"2b",
          3667 => x"06",
          3668 => x"51",
          3669 => x"53",
          3670 => x"88",
          3671 => x"72",
          3672 => x"74",
          3673 => x"82",
          3674 => x"70",
          3675 => x"81",
          3676 => x"8b",
          3677 => x"2b",
          3678 => x"57",
          3679 => x"70",
          3680 => x"33",
          3681 => x"07",
          3682 => x"ff",
          3683 => x"2a",
          3684 => x"58",
          3685 => x"34",
          3686 => x"34",
          3687 => x"04",
          3688 => x"82",
          3689 => x"02",
          3690 => x"05",
          3691 => x"2b",
          3692 => x"11",
          3693 => x"33",
          3694 => x"71",
          3695 => x"59",
          3696 => x"56",
          3697 => x"71",
          3698 => x"33",
          3699 => x"07",
          3700 => x"a2",
          3701 => x"07",
          3702 => x"53",
          3703 => x"53",
          3704 => x"70",
          3705 => x"82",
          3706 => x"70",
          3707 => x"81",
          3708 => x"8b",
          3709 => x"2b",
          3710 => x"57",
          3711 => x"82",
          3712 => x"13",
          3713 => x"2b",
          3714 => x"2a",
          3715 => x"52",
          3716 => x"34",
          3717 => x"34",
          3718 => x"08",
          3719 => x"33",
          3720 => x"71",
          3721 => x"82",
          3722 => x"52",
          3723 => x"0d",
          3724 => x"0d",
          3725 => x"e4",
          3726 => x"2a",
          3727 => x"ff",
          3728 => x"57",
          3729 => x"3f",
          3730 => x"08",
          3731 => x"71",
          3732 => x"33",
          3733 => x"71",
          3734 => x"83",
          3735 => x"11",
          3736 => x"12",
          3737 => x"2b",
          3738 => x"07",
          3739 => x"51",
          3740 => x"55",
          3741 => x"80",
          3742 => x"82",
          3743 => x"75",
          3744 => x"3f",
          3745 => x"84",
          3746 => x"15",
          3747 => x"2b",
          3748 => x"07",
          3749 => x"88",
          3750 => x"55",
          3751 => x"86",
          3752 => x"81",
          3753 => x"75",
          3754 => x"82",
          3755 => x"70",
          3756 => x"33",
          3757 => x"71",
          3758 => x"70",
          3759 => x"57",
          3760 => x"72",
          3761 => x"73",
          3762 => x"82",
          3763 => x"18",
          3764 => x"86",
          3765 => x"0b",
          3766 => x"82",
          3767 => x"53",
          3768 => x"34",
          3769 => x"34",
          3770 => x"08",
          3771 => x"81",
          3772 => x"88",
          3773 => x"82",
          3774 => x"70",
          3775 => x"51",
          3776 => x"74",
          3777 => x"81",
          3778 => x"3d",
          3779 => x"3d",
          3780 => x"82",
          3781 => x"84",
          3782 => x"3f",
          3783 => x"86",
          3784 => x"fe",
          3785 => x"3d",
          3786 => x"3d",
          3787 => x"52",
          3788 => x"3f",
          3789 => x"08",
          3790 => x"06",
          3791 => x"08",
          3792 => x"85",
          3793 => x"88",
          3794 => x"5f",
          3795 => x"5a",
          3796 => x"59",
          3797 => x"80",
          3798 => x"83",
          3799 => x"70",
          3800 => x"33",
          3801 => x"07",
          3802 => x"ff",
          3803 => x"70",
          3804 => x"06",
          3805 => x"52",
          3806 => x"59",
          3807 => x"27",
          3808 => x"80",
          3809 => x"75",
          3810 => x"84",
          3811 => x"16",
          3812 => x"2b",
          3813 => x"75",
          3814 => x"81",
          3815 => x"85",
          3816 => x"59",
          3817 => x"83",
          3818 => x"e4",
          3819 => x"33",
          3820 => x"71",
          3821 => x"70",
          3822 => x"06",
          3823 => x"56",
          3824 => x"75",
          3825 => x"81",
          3826 => x"79",
          3827 => x"cc",
          3828 => x"74",
          3829 => x"c4",
          3830 => x"2e",
          3831 => x"89",
          3832 => x"f8",
          3833 => x"ac",
          3834 => x"80",
          3835 => x"75",
          3836 => x"3f",
          3837 => x"08",
          3838 => x"11",
          3839 => x"33",
          3840 => x"71",
          3841 => x"53",
          3842 => x"74",
          3843 => x"70",
          3844 => x"06",
          3845 => x"5c",
          3846 => x"78",
          3847 => x"76",
          3848 => x"57",
          3849 => x"34",
          3850 => x"08",
          3851 => x"71",
          3852 => x"86",
          3853 => x"12",
          3854 => x"2b",
          3855 => x"2a",
          3856 => x"53",
          3857 => x"73",
          3858 => x"75",
          3859 => x"82",
          3860 => x"70",
          3861 => x"33",
          3862 => x"71",
          3863 => x"83",
          3864 => x"5d",
          3865 => x"05",
          3866 => x"15",
          3867 => x"15",
          3868 => x"e4",
          3869 => x"71",
          3870 => x"33",
          3871 => x"71",
          3872 => x"70",
          3873 => x"5a",
          3874 => x"54",
          3875 => x"34",
          3876 => x"34",
          3877 => x"08",
          3878 => x"54",
          3879 => x"ec",
          3880 => x"0d",
          3881 => x"0d",
          3882 => x"85",
          3883 => x"38",
          3884 => x"71",
          3885 => x"2e",
          3886 => x"51",
          3887 => x"82",
          3888 => x"53",
          3889 => x"ec",
          3890 => x"0d",
          3891 => x"0d",
          3892 => x"33",
          3893 => x"70",
          3894 => x"38",
          3895 => x"11",
          3896 => x"82",
          3897 => x"83",
          3898 => x"fc",
          3899 => x"9b",
          3900 => x"84",
          3901 => x"33",
          3902 => x"51",
          3903 => x"80",
          3904 => x"84",
          3905 => x"92",
          3906 => x"51",
          3907 => x"80",
          3908 => x"81",
          3909 => x"72",
          3910 => x"92",
          3911 => x"81",
          3912 => x"0b",
          3913 => x"8c",
          3914 => x"71",
          3915 => x"06",
          3916 => x"80",
          3917 => x"87",
          3918 => x"08",
          3919 => x"38",
          3920 => x"80",
          3921 => x"71",
          3922 => x"c0",
          3923 => x"51",
          3924 => x"87",
          3925 => x"85",
          3926 => x"82",
          3927 => x"33",
          3928 => x"85",
          3929 => x"3d",
          3930 => x"3d",
          3931 => x"64",
          3932 => x"bf",
          3933 => x"40",
          3934 => x"74",
          3935 => x"cd",
          3936 => x"ec",
          3937 => x"7a",
          3938 => x"81",
          3939 => x"72",
          3940 => x"87",
          3941 => x"11",
          3942 => x"8c",
          3943 => x"92",
          3944 => x"5a",
          3945 => x"58",
          3946 => x"c0",
          3947 => x"76",
          3948 => x"76",
          3949 => x"70",
          3950 => x"81",
          3951 => x"54",
          3952 => x"8e",
          3953 => x"52",
          3954 => x"81",
          3955 => x"81",
          3956 => x"74",
          3957 => x"53",
          3958 => x"83",
          3959 => x"78",
          3960 => x"8f",
          3961 => x"2e",
          3962 => x"c0",
          3963 => x"52",
          3964 => x"87",
          3965 => x"08",
          3966 => x"2e",
          3967 => x"84",
          3968 => x"38",
          3969 => x"87",
          3970 => x"15",
          3971 => x"70",
          3972 => x"52",
          3973 => x"ff",
          3974 => x"39",
          3975 => x"81",
          3976 => x"ff",
          3977 => x"57",
          3978 => x"90",
          3979 => x"80",
          3980 => x"71",
          3981 => x"78",
          3982 => x"38",
          3983 => x"80",
          3984 => x"80",
          3985 => x"81",
          3986 => x"72",
          3987 => x"0c",
          3988 => x"04",
          3989 => x"60",
          3990 => x"8c",
          3991 => x"33",
          3992 => x"5b",
          3993 => x"74",
          3994 => x"e1",
          3995 => x"ec",
          3996 => x"79",
          3997 => x"78",
          3998 => x"06",
          3999 => x"77",
          4000 => x"87",
          4001 => x"11",
          4002 => x"8c",
          4003 => x"92",
          4004 => x"59",
          4005 => x"85",
          4006 => x"98",
          4007 => x"7d",
          4008 => x"0c",
          4009 => x"08",
          4010 => x"70",
          4011 => x"53",
          4012 => x"2e",
          4013 => x"70",
          4014 => x"33",
          4015 => x"18",
          4016 => x"2a",
          4017 => x"51",
          4018 => x"2e",
          4019 => x"c0",
          4020 => x"52",
          4021 => x"87",
          4022 => x"08",
          4023 => x"2e",
          4024 => x"84",
          4025 => x"38",
          4026 => x"87",
          4027 => x"15",
          4028 => x"70",
          4029 => x"52",
          4030 => x"ff",
          4031 => x"39",
          4032 => x"81",
          4033 => x"80",
          4034 => x"52",
          4035 => x"90",
          4036 => x"80",
          4037 => x"71",
          4038 => x"7a",
          4039 => x"38",
          4040 => x"80",
          4041 => x"80",
          4042 => x"81",
          4043 => x"72",
          4044 => x"0c",
          4045 => x"04",
          4046 => x"7a",
          4047 => x"a3",
          4048 => x"88",
          4049 => x"33",
          4050 => x"56",
          4051 => x"3f",
          4052 => x"08",
          4053 => x"83",
          4054 => x"fe",
          4055 => x"87",
          4056 => x"0c",
          4057 => x"76",
          4058 => x"38",
          4059 => x"93",
          4060 => x"2b",
          4061 => x"8c",
          4062 => x"71",
          4063 => x"38",
          4064 => x"71",
          4065 => x"c6",
          4066 => x"39",
          4067 => x"81",
          4068 => x"06",
          4069 => x"71",
          4070 => x"38",
          4071 => x"8c",
          4072 => x"e8",
          4073 => x"98",
          4074 => x"71",
          4075 => x"73",
          4076 => x"92",
          4077 => x"72",
          4078 => x"06",
          4079 => x"f7",
          4080 => x"80",
          4081 => x"88",
          4082 => x"0c",
          4083 => x"80",
          4084 => x"56",
          4085 => x"56",
          4086 => x"82",
          4087 => x"88",
          4088 => x"fe",
          4089 => x"81",
          4090 => x"33",
          4091 => x"07",
          4092 => x"0c",
          4093 => x"3d",
          4094 => x"3d",
          4095 => x"11",
          4096 => x"33",
          4097 => x"71",
          4098 => x"81",
          4099 => x"72",
          4100 => x"75",
          4101 => x"82",
          4102 => x"52",
          4103 => x"54",
          4104 => x"0d",
          4105 => x"0d",
          4106 => x"05",
          4107 => x"52",
          4108 => x"70",
          4109 => x"34",
          4110 => x"51",
          4111 => x"83",
          4112 => x"ff",
          4113 => x"75",
          4114 => x"72",
          4115 => x"54",
          4116 => x"2a",
          4117 => x"70",
          4118 => x"34",
          4119 => x"51",
          4120 => x"81",
          4121 => x"70",
          4122 => x"70",
          4123 => x"3d",
          4124 => x"3d",
          4125 => x"77",
          4126 => x"70",
          4127 => x"38",
          4128 => x"05",
          4129 => x"70",
          4130 => x"34",
          4131 => x"eb",
          4132 => x"0d",
          4133 => x"0d",
          4134 => x"54",
          4135 => x"72",
          4136 => x"54",
          4137 => x"51",
          4138 => x"84",
          4139 => x"fc",
          4140 => x"77",
          4141 => x"53",
          4142 => x"05",
          4143 => x"70",
          4144 => x"33",
          4145 => x"ff",
          4146 => x"52",
          4147 => x"2e",
          4148 => x"80",
          4149 => x"71",
          4150 => x"0c",
          4151 => x"04",
          4152 => x"74",
          4153 => x"89",
          4154 => x"2e",
          4155 => x"11",
          4156 => x"52",
          4157 => x"70",
          4158 => x"ec",
          4159 => x"0d",
          4160 => x"82",
          4161 => x"04",
          4162 => x"85",
          4163 => x"f7",
          4164 => x"56",
          4165 => x"17",
          4166 => x"74",
          4167 => x"d6",
          4168 => x"b0",
          4169 => x"b4",
          4170 => x"81",
          4171 => x"59",
          4172 => x"82",
          4173 => x"7a",
          4174 => x"06",
          4175 => x"85",
          4176 => x"17",
          4177 => x"08",
          4178 => x"08",
          4179 => x"08",
          4180 => x"74",
          4181 => x"38",
          4182 => x"55",
          4183 => x"09",
          4184 => x"38",
          4185 => x"18",
          4186 => x"81",
          4187 => x"f9",
          4188 => x"39",
          4189 => x"82",
          4190 => x"8b",
          4191 => x"fa",
          4192 => x"7a",
          4193 => x"57",
          4194 => x"08",
          4195 => x"75",
          4196 => x"3f",
          4197 => x"08",
          4198 => x"ec",
          4199 => x"81",
          4200 => x"b4",
          4201 => x"16",
          4202 => x"be",
          4203 => x"ec",
          4204 => x"85",
          4205 => x"81",
          4206 => x"17",
          4207 => x"85",
          4208 => x"3d",
          4209 => x"3d",
          4210 => x"52",
          4211 => x"3f",
          4212 => x"08",
          4213 => x"ec",
          4214 => x"38",
          4215 => x"74",
          4216 => x"81",
          4217 => x"38",
          4218 => x"59",
          4219 => x"09",
          4220 => x"e3",
          4221 => x"53",
          4222 => x"08",
          4223 => x"70",
          4224 => x"91",
          4225 => x"d5",
          4226 => x"17",
          4227 => x"3f",
          4228 => x"a4",
          4229 => x"51",
          4230 => x"86",
          4231 => x"f2",
          4232 => x"17",
          4233 => x"3f",
          4234 => x"52",
          4235 => x"51",
          4236 => x"8c",
          4237 => x"84",
          4238 => x"fc",
          4239 => x"17",
          4240 => x"70",
          4241 => x"79",
          4242 => x"52",
          4243 => x"51",
          4244 => x"77",
          4245 => x"80",
          4246 => x"81",
          4247 => x"f9",
          4248 => x"85",
          4249 => x"2e",
          4250 => x"58",
          4251 => x"ec",
          4252 => x"0d",
          4253 => x"0d",
          4254 => x"98",
          4255 => x"05",
          4256 => x"80",
          4257 => x"27",
          4258 => x"15",
          4259 => x"51",
          4260 => x"3f",
          4261 => x"82",
          4262 => x"05",
          4263 => x"85",
          4264 => x"3d",
          4265 => x"3d",
          4266 => x"70",
          4267 => x"57",
          4268 => x"81",
          4269 => x"98",
          4270 => x"81",
          4271 => x"74",
          4272 => x"72",
          4273 => x"f5",
          4274 => x"24",
          4275 => x"81",
          4276 => x"81",
          4277 => x"83",
          4278 => x"38",
          4279 => x"76",
          4280 => x"70",
          4281 => x"16",
          4282 => x"74",
          4283 => x"8f",
          4284 => x"ec",
          4285 => x"38",
          4286 => x"06",
          4287 => x"33",
          4288 => x"89",
          4289 => x"08",
          4290 => x"54",
          4291 => x"fc",
          4292 => x"85",
          4293 => x"fe",
          4294 => x"ff",
          4295 => x"11",
          4296 => x"2b",
          4297 => x"81",
          4298 => x"2a",
          4299 => x"51",
          4300 => x"e2",
          4301 => x"ff",
          4302 => x"da",
          4303 => x"2a",
          4304 => x"05",
          4305 => x"fc",
          4306 => x"85",
          4307 => x"c6",
          4308 => x"83",
          4309 => x"05",
          4310 => x"f9",
          4311 => x"85",
          4312 => x"ff",
          4313 => x"ae",
          4314 => x"2a",
          4315 => x"05",
          4316 => x"fc",
          4317 => x"85",
          4318 => x"38",
          4319 => x"83",
          4320 => x"05",
          4321 => x"f8",
          4322 => x"85",
          4323 => x"0a",
          4324 => x"39",
          4325 => x"82",
          4326 => x"89",
          4327 => x"f8",
          4328 => x"7c",
          4329 => x"56",
          4330 => x"77",
          4331 => x"38",
          4332 => x"08",
          4333 => x"38",
          4334 => x"72",
          4335 => x"9d",
          4336 => x"24",
          4337 => x"81",
          4338 => x"82",
          4339 => x"83",
          4340 => x"38",
          4341 => x"76",
          4342 => x"70",
          4343 => x"18",
          4344 => x"76",
          4345 => x"97",
          4346 => x"ec",
          4347 => x"85",
          4348 => x"d9",
          4349 => x"ff",
          4350 => x"05",
          4351 => x"81",
          4352 => x"54",
          4353 => x"80",
          4354 => x"77",
          4355 => x"f0",
          4356 => x"8f",
          4357 => x"51",
          4358 => x"34",
          4359 => x"17",
          4360 => x"2a",
          4361 => x"05",
          4362 => x"fa",
          4363 => x"85",
          4364 => x"82",
          4365 => x"81",
          4366 => x"83",
          4367 => x"b4",
          4368 => x"2a",
          4369 => x"8f",
          4370 => x"2a",
          4371 => x"f0",
          4372 => x"06",
          4373 => x"72",
          4374 => x"ec",
          4375 => x"2a",
          4376 => x"05",
          4377 => x"fa",
          4378 => x"85",
          4379 => x"82",
          4380 => x"80",
          4381 => x"83",
          4382 => x"52",
          4383 => x"fe",
          4384 => x"b4",
          4385 => x"9d",
          4386 => x"76",
          4387 => x"17",
          4388 => x"75",
          4389 => x"3f",
          4390 => x"08",
          4391 => x"ec",
          4392 => x"77",
          4393 => x"77",
          4394 => x"fc",
          4395 => x"b4",
          4396 => x"51",
          4397 => x"c2",
          4398 => x"ec",
          4399 => x"06",
          4400 => x"72",
          4401 => x"3f",
          4402 => x"17",
          4403 => x"85",
          4404 => x"3d",
          4405 => x"3d",
          4406 => x"7e",
          4407 => x"56",
          4408 => x"75",
          4409 => x"74",
          4410 => x"27",
          4411 => x"80",
          4412 => x"ff",
          4413 => x"75",
          4414 => x"3f",
          4415 => x"08",
          4416 => x"ec",
          4417 => x"38",
          4418 => x"54",
          4419 => x"81",
          4420 => x"39",
          4421 => x"08",
          4422 => x"39",
          4423 => x"51",
          4424 => x"82",
          4425 => x"58",
          4426 => x"08",
          4427 => x"c7",
          4428 => x"ec",
          4429 => x"d2",
          4430 => x"ec",
          4431 => x"cf",
          4432 => x"74",
          4433 => x"fc",
          4434 => x"85",
          4435 => x"38",
          4436 => x"fe",
          4437 => x"08",
          4438 => x"74",
          4439 => x"38",
          4440 => x"17",
          4441 => x"33",
          4442 => x"73",
          4443 => x"77",
          4444 => x"26",
          4445 => x"80",
          4446 => x"85",
          4447 => x"3d",
          4448 => x"3d",
          4449 => x"71",
          4450 => x"5b",
          4451 => x"8c",
          4452 => x"77",
          4453 => x"38",
          4454 => x"78",
          4455 => x"81",
          4456 => x"79",
          4457 => x"f9",
          4458 => x"55",
          4459 => x"ec",
          4460 => x"e6",
          4461 => x"ec",
          4462 => x"85",
          4463 => x"2e",
          4464 => x"98",
          4465 => x"85",
          4466 => x"82",
          4467 => x"58",
          4468 => x"70",
          4469 => x"80",
          4470 => x"38",
          4471 => x"09",
          4472 => x"e4",
          4473 => x"56",
          4474 => x"76",
          4475 => x"82",
          4476 => x"7a",
          4477 => x"3f",
          4478 => x"85",
          4479 => x"2e",
          4480 => x"86",
          4481 => x"ec",
          4482 => x"85",
          4483 => x"70",
          4484 => x"70",
          4485 => x"25",
          4486 => x"82",
          4487 => x"54",
          4488 => x"55",
          4489 => x"38",
          4490 => x"08",
          4491 => x"38",
          4492 => x"54",
          4493 => x"90",
          4494 => x"18",
          4495 => x"38",
          4496 => x"39",
          4497 => x"38",
          4498 => x"16",
          4499 => x"08",
          4500 => x"38",
          4501 => x"78",
          4502 => x"38",
          4503 => x"51",
          4504 => x"82",
          4505 => x"80",
          4506 => x"80",
          4507 => x"ec",
          4508 => x"09",
          4509 => x"38",
          4510 => x"08",
          4511 => x"ec",
          4512 => x"09",
          4513 => x"72",
          4514 => x"70",
          4515 => x"51",
          4516 => x"80",
          4517 => x"78",
          4518 => x"06",
          4519 => x"73",
          4520 => x"39",
          4521 => x"52",
          4522 => x"f3",
          4523 => x"ec",
          4524 => x"ec",
          4525 => x"05",
          4526 => x"ec",
          4527 => x"25",
          4528 => x"79",
          4529 => x"38",
          4530 => x"8f",
          4531 => x"79",
          4532 => x"f9",
          4533 => x"85",
          4534 => x"74",
          4535 => x"8c",
          4536 => x"17",
          4537 => x"90",
          4538 => x"54",
          4539 => x"86",
          4540 => x"90",
          4541 => x"17",
          4542 => x"54",
          4543 => x"34",
          4544 => x"56",
          4545 => x"90",
          4546 => x"80",
          4547 => x"82",
          4548 => x"55",
          4549 => x"56",
          4550 => x"82",
          4551 => x"8c",
          4552 => x"f8",
          4553 => x"70",
          4554 => x"e3",
          4555 => x"ec",
          4556 => x"56",
          4557 => x"08",
          4558 => x"7b",
          4559 => x"f6",
          4560 => x"85",
          4561 => x"85",
          4562 => x"17",
          4563 => x"80",
          4564 => x"b4",
          4565 => x"57",
          4566 => x"77",
          4567 => x"81",
          4568 => x"15",
          4569 => x"78",
          4570 => x"81",
          4571 => x"53",
          4572 => x"15",
          4573 => x"dc",
          4574 => x"ec",
          4575 => x"df",
          4576 => x"22",
          4577 => x"09",
          4578 => x"72",
          4579 => x"2a",
          4580 => x"56",
          4581 => x"ec",
          4582 => x"0d",
          4583 => x"0d",
          4584 => x"08",
          4585 => x"74",
          4586 => x"26",
          4587 => x"74",
          4588 => x"72",
          4589 => x"74",
          4590 => x"88",
          4591 => x"73",
          4592 => x"33",
          4593 => x"27",
          4594 => x"16",
          4595 => x"9b",
          4596 => x"2a",
          4597 => x"88",
          4598 => x"58",
          4599 => x"80",
          4600 => x"16",
          4601 => x"0c",
          4602 => x"8a",
          4603 => x"89",
          4604 => x"72",
          4605 => x"38",
          4606 => x"51",
          4607 => x"82",
          4608 => x"54",
          4609 => x"08",
          4610 => x"38",
          4611 => x"85",
          4612 => x"8b",
          4613 => x"08",
          4614 => x"08",
          4615 => x"82",
          4616 => x"74",
          4617 => x"cb",
          4618 => x"75",
          4619 => x"3f",
          4620 => x"08",
          4621 => x"73",
          4622 => x"98",
          4623 => x"82",
          4624 => x"2e",
          4625 => x"39",
          4626 => x"39",
          4627 => x"13",
          4628 => x"74",
          4629 => x"16",
          4630 => x"18",
          4631 => x"77",
          4632 => x"0c",
          4633 => x"04",
          4634 => x"7a",
          4635 => x"12",
          4636 => x"59",
          4637 => x"80",
          4638 => x"86",
          4639 => x"98",
          4640 => x"14",
          4641 => x"55",
          4642 => x"81",
          4643 => x"83",
          4644 => x"77",
          4645 => x"81",
          4646 => x"0c",
          4647 => x"55",
          4648 => x"76",
          4649 => x"17",
          4650 => x"74",
          4651 => x"9b",
          4652 => x"39",
          4653 => x"ff",
          4654 => x"2a",
          4655 => x"81",
          4656 => x"52",
          4657 => x"de",
          4658 => x"ec",
          4659 => x"55",
          4660 => x"85",
          4661 => x"80",
          4662 => x"55",
          4663 => x"08",
          4664 => x"f4",
          4665 => x"08",
          4666 => x"08",
          4667 => x"38",
          4668 => x"77",
          4669 => x"84",
          4670 => x"39",
          4671 => x"52",
          4672 => x"fe",
          4673 => x"ec",
          4674 => x"55",
          4675 => x"08",
          4676 => x"c4",
          4677 => x"82",
          4678 => x"81",
          4679 => x"81",
          4680 => x"ec",
          4681 => x"b0",
          4682 => x"ec",
          4683 => x"51",
          4684 => x"82",
          4685 => x"a0",
          4686 => x"15",
          4687 => x"75",
          4688 => x"3f",
          4689 => x"08",
          4690 => x"76",
          4691 => x"77",
          4692 => x"9c",
          4693 => x"55",
          4694 => x"ec",
          4695 => x"0d",
          4696 => x"0d",
          4697 => x"08",
          4698 => x"80",
          4699 => x"fc",
          4700 => x"85",
          4701 => x"82",
          4702 => x"80",
          4703 => x"85",
          4704 => x"98",
          4705 => x"78",
          4706 => x"3f",
          4707 => x"08",
          4708 => x"ec",
          4709 => x"38",
          4710 => x"08",
          4711 => x"70",
          4712 => x"58",
          4713 => x"2e",
          4714 => x"83",
          4715 => x"82",
          4716 => x"55",
          4717 => x"81",
          4718 => x"07",
          4719 => x"2e",
          4720 => x"16",
          4721 => x"2e",
          4722 => x"88",
          4723 => x"82",
          4724 => x"56",
          4725 => x"51",
          4726 => x"82",
          4727 => x"54",
          4728 => x"08",
          4729 => x"9b",
          4730 => x"2e",
          4731 => x"83",
          4732 => x"73",
          4733 => x"0c",
          4734 => x"04",
          4735 => x"76",
          4736 => x"54",
          4737 => x"82",
          4738 => x"83",
          4739 => x"76",
          4740 => x"53",
          4741 => x"2e",
          4742 => x"90",
          4743 => x"51",
          4744 => x"82",
          4745 => x"90",
          4746 => x"53",
          4747 => x"ec",
          4748 => x"0d",
          4749 => x"0d",
          4750 => x"83",
          4751 => x"54",
          4752 => x"55",
          4753 => x"3f",
          4754 => x"51",
          4755 => x"2e",
          4756 => x"8b",
          4757 => x"2a",
          4758 => x"51",
          4759 => x"86",
          4760 => x"f7",
          4761 => x"7d",
          4762 => x"75",
          4763 => x"98",
          4764 => x"2e",
          4765 => x"98",
          4766 => x"78",
          4767 => x"3f",
          4768 => x"08",
          4769 => x"ec",
          4770 => x"38",
          4771 => x"70",
          4772 => x"73",
          4773 => x"58",
          4774 => x"8b",
          4775 => x"bf",
          4776 => x"ff",
          4777 => x"53",
          4778 => x"34",
          4779 => x"08",
          4780 => x"e5",
          4781 => x"81",
          4782 => x"2e",
          4783 => x"70",
          4784 => x"57",
          4785 => x"9e",
          4786 => x"2e",
          4787 => x"85",
          4788 => x"df",
          4789 => x"72",
          4790 => x"81",
          4791 => x"76",
          4792 => x"2e",
          4793 => x"52",
          4794 => x"fc",
          4795 => x"ec",
          4796 => x"85",
          4797 => x"38",
          4798 => x"fe",
          4799 => x"39",
          4800 => x"16",
          4801 => x"85",
          4802 => x"3d",
          4803 => x"3d",
          4804 => x"08",
          4805 => x"52",
          4806 => x"c5",
          4807 => x"ec",
          4808 => x"85",
          4809 => x"38",
          4810 => x"52",
          4811 => x"cf",
          4812 => x"ec",
          4813 => x"85",
          4814 => x"38",
          4815 => x"85",
          4816 => x"9c",
          4817 => x"ea",
          4818 => x"53",
          4819 => x"9c",
          4820 => x"ea",
          4821 => x"0b",
          4822 => x"74",
          4823 => x"0c",
          4824 => x"04",
          4825 => x"75",
          4826 => x"12",
          4827 => x"53",
          4828 => x"8b",
          4829 => x"ec",
          4830 => x"9c",
          4831 => x"e5",
          4832 => x"0b",
          4833 => x"85",
          4834 => x"fa",
          4835 => x"7a",
          4836 => x"0b",
          4837 => x"98",
          4838 => x"2e",
          4839 => x"80",
          4840 => x"55",
          4841 => x"17",
          4842 => x"33",
          4843 => x"51",
          4844 => x"2e",
          4845 => x"85",
          4846 => x"06",
          4847 => x"e5",
          4848 => x"2e",
          4849 => x"8b",
          4850 => x"70",
          4851 => x"34",
          4852 => x"71",
          4853 => x"05",
          4854 => x"15",
          4855 => x"27",
          4856 => x"15",
          4857 => x"80",
          4858 => x"34",
          4859 => x"52",
          4860 => x"88",
          4861 => x"17",
          4862 => x"52",
          4863 => x"3f",
          4864 => x"08",
          4865 => x"12",
          4866 => x"3f",
          4867 => x"08",
          4868 => x"98",
          4869 => x"cb",
          4870 => x"ec",
          4871 => x"23",
          4872 => x"04",
          4873 => x"7f",
          4874 => x"5b",
          4875 => x"33",
          4876 => x"73",
          4877 => x"38",
          4878 => x"80",
          4879 => x"38",
          4880 => x"8c",
          4881 => x"08",
          4882 => x"ac",
          4883 => x"41",
          4884 => x"33",
          4885 => x"73",
          4886 => x"81",
          4887 => x"81",
          4888 => x"dc",
          4889 => x"81",
          4890 => x"25",
          4891 => x"51",
          4892 => x"38",
          4893 => x"0c",
          4894 => x"51",
          4895 => x"26",
          4896 => x"80",
          4897 => x"34",
          4898 => x"51",
          4899 => x"82",
          4900 => x"55",
          4901 => x"91",
          4902 => x"1d",
          4903 => x"8b",
          4904 => x"79",
          4905 => x"3f",
          4906 => x"57",
          4907 => x"55",
          4908 => x"2e",
          4909 => x"80",
          4910 => x"18",
          4911 => x"1a",
          4912 => x"70",
          4913 => x"70",
          4914 => x"82",
          4915 => x"51",
          4916 => x"54",
          4917 => x"79",
          4918 => x"74",
          4919 => x"57",
          4920 => x"af",
          4921 => x"81",
          4922 => x"2a",
          4923 => x"75",
          4924 => x"8c",
          4925 => x"2e",
          4926 => x"a0",
          4927 => x"38",
          4928 => x"0c",
          4929 => x"76",
          4930 => x"38",
          4931 => x"c2",
          4932 => x"70",
          4933 => x"5a",
          4934 => x"76",
          4935 => x"38",
          4936 => x"70",
          4937 => x"77",
          4938 => x"70",
          4939 => x"72",
          4940 => x"80",
          4941 => x"51",
          4942 => x"73",
          4943 => x"38",
          4944 => x"18",
          4945 => x"1a",
          4946 => x"55",
          4947 => x"2e",
          4948 => x"83",
          4949 => x"73",
          4950 => x"70",
          4951 => x"70",
          4952 => x"07",
          4953 => x"73",
          4954 => x"b9",
          4955 => x"2e",
          4956 => x"83",
          4957 => x"76",
          4958 => x"07",
          4959 => x"2e",
          4960 => x"8b",
          4961 => x"81",
          4962 => x"32",
          4963 => x"05",
          4964 => x"71",
          4965 => x"53",
          4966 => x"55",
          4967 => x"38",
          4968 => x"5c",
          4969 => x"75",
          4970 => x"73",
          4971 => x"38",
          4972 => x"06",
          4973 => x"11",
          4974 => x"75",
          4975 => x"3f",
          4976 => x"08",
          4977 => x"38",
          4978 => x"33",
          4979 => x"54",
          4980 => x"e6",
          4981 => x"85",
          4982 => x"2e",
          4983 => x"ff",
          4984 => x"74",
          4985 => x"38",
          4986 => x"75",
          4987 => x"17",
          4988 => x"57",
          4989 => x"a7",
          4990 => x"81",
          4991 => x"e5",
          4992 => x"85",
          4993 => x"38",
          4994 => x"54",
          4995 => x"89",
          4996 => x"70",
          4997 => x"57",
          4998 => x"54",
          4999 => x"81",
          5000 => x"ed",
          5001 => x"7e",
          5002 => x"2e",
          5003 => x"33",
          5004 => x"e5",
          5005 => x"06",
          5006 => x"7a",
          5007 => x"a0",
          5008 => x"38",
          5009 => x"55",
          5010 => x"84",
          5011 => x"39",
          5012 => x"8b",
          5013 => x"7b",
          5014 => x"7a",
          5015 => x"3f",
          5016 => x"08",
          5017 => x"ec",
          5018 => x"38",
          5019 => x"52",
          5020 => x"8b",
          5021 => x"ec",
          5022 => x"85",
          5023 => x"c2",
          5024 => x"08",
          5025 => x"55",
          5026 => x"ff",
          5027 => x"15",
          5028 => x"54",
          5029 => x"34",
          5030 => x"70",
          5031 => x"81",
          5032 => x"58",
          5033 => x"8b",
          5034 => x"74",
          5035 => x"3f",
          5036 => x"08",
          5037 => x"38",
          5038 => x"51",
          5039 => x"ff",
          5040 => x"ab",
          5041 => x"55",
          5042 => x"bb",
          5043 => x"2e",
          5044 => x"80",
          5045 => x"85",
          5046 => x"06",
          5047 => x"58",
          5048 => x"80",
          5049 => x"75",
          5050 => x"73",
          5051 => x"a7",
          5052 => x"0b",
          5053 => x"80",
          5054 => x"39",
          5055 => x"54",
          5056 => x"85",
          5057 => x"75",
          5058 => x"81",
          5059 => x"73",
          5060 => x"1b",
          5061 => x"2a",
          5062 => x"51",
          5063 => x"80",
          5064 => x"90",
          5065 => x"ff",
          5066 => x"05",
          5067 => x"f5",
          5068 => x"85",
          5069 => x"1c",
          5070 => x"39",
          5071 => x"ec",
          5072 => x"0d",
          5073 => x"0d",
          5074 => x"7b",
          5075 => x"73",
          5076 => x"55",
          5077 => x"2e",
          5078 => x"75",
          5079 => x"57",
          5080 => x"26",
          5081 => x"ba",
          5082 => x"70",
          5083 => x"ba",
          5084 => x"06",
          5085 => x"73",
          5086 => x"70",
          5087 => x"51",
          5088 => x"89",
          5089 => x"82",
          5090 => x"ff",
          5091 => x"56",
          5092 => x"2e",
          5093 => x"80",
          5094 => x"a4",
          5095 => x"08",
          5096 => x"76",
          5097 => x"58",
          5098 => x"81",
          5099 => x"ff",
          5100 => x"53",
          5101 => x"26",
          5102 => x"13",
          5103 => x"06",
          5104 => x"9f",
          5105 => x"99",
          5106 => x"e0",
          5107 => x"ff",
          5108 => x"72",
          5109 => x"70",
          5110 => x"51",
          5111 => x"09",
          5112 => x"38",
          5113 => x"38",
          5114 => x"05",
          5115 => x"70",
          5116 => x"70",
          5117 => x"2a",
          5118 => x"07",
          5119 => x"51",
          5120 => x"8f",
          5121 => x"84",
          5122 => x"83",
          5123 => x"8e",
          5124 => x"74",
          5125 => x"38",
          5126 => x"0c",
          5127 => x"86",
          5128 => x"a4",
          5129 => x"82",
          5130 => x"8c",
          5131 => x"fa",
          5132 => x"56",
          5133 => x"17",
          5134 => x"b0",
          5135 => x"52",
          5136 => x"bb",
          5137 => x"82",
          5138 => x"81",
          5139 => x"b2",
          5140 => x"8f",
          5141 => x"ec",
          5142 => x"ff",
          5143 => x"55",
          5144 => x"d5",
          5145 => x"06",
          5146 => x"80",
          5147 => x"33",
          5148 => x"81",
          5149 => x"81",
          5150 => x"81",
          5151 => x"eb",
          5152 => x"81",
          5153 => x"25",
          5154 => x"51",
          5155 => x"38",
          5156 => x"2e",
          5157 => x"b5",
          5158 => x"81",
          5159 => x"80",
          5160 => x"e0",
          5161 => x"85",
          5162 => x"82",
          5163 => x"80",
          5164 => x"85",
          5165 => x"e8",
          5166 => x"16",
          5167 => x"3f",
          5168 => x"08",
          5169 => x"ec",
          5170 => x"83",
          5171 => x"74",
          5172 => x"0c",
          5173 => x"04",
          5174 => x"62",
          5175 => x"80",
          5176 => x"58",
          5177 => x"0c",
          5178 => x"d9",
          5179 => x"ec",
          5180 => x"56",
          5181 => x"85",
          5182 => x"87",
          5183 => x"85",
          5184 => x"2b",
          5185 => x"11",
          5186 => x"8c",
          5187 => x"2e",
          5188 => x"73",
          5189 => x"81",
          5190 => x"33",
          5191 => x"80",
          5192 => x"81",
          5193 => x"d7",
          5194 => x"85",
          5195 => x"ff",
          5196 => x"06",
          5197 => x"98",
          5198 => x"2e",
          5199 => x"74",
          5200 => x"81",
          5201 => x"8a",
          5202 => x"b4",
          5203 => x"39",
          5204 => x"77",
          5205 => x"81",
          5206 => x"33",
          5207 => x"3f",
          5208 => x"08",
          5209 => x"70",
          5210 => x"55",
          5211 => x"86",
          5212 => x"80",
          5213 => x"74",
          5214 => x"81",
          5215 => x"8a",
          5216 => x"fc",
          5217 => x"53",
          5218 => x"fd",
          5219 => x"85",
          5220 => x"ff",
          5221 => x"82",
          5222 => x"06",
          5223 => x"8d",
          5224 => x"58",
          5225 => x"f6",
          5226 => x"58",
          5227 => x"2e",
          5228 => x"fa",
          5229 => x"c2",
          5230 => x"ec",
          5231 => x"78",
          5232 => x"5a",
          5233 => x"90",
          5234 => x"75",
          5235 => x"38",
          5236 => x"3d",
          5237 => x"70",
          5238 => x"08",
          5239 => x"7b",
          5240 => x"38",
          5241 => x"51",
          5242 => x"82",
          5243 => x"81",
          5244 => x"81",
          5245 => x"38",
          5246 => x"83",
          5247 => x"38",
          5248 => x"84",
          5249 => x"38",
          5250 => x"81",
          5251 => x"38",
          5252 => x"db",
          5253 => x"85",
          5254 => x"ff",
          5255 => x"72",
          5256 => x"09",
          5257 => x"d8",
          5258 => x"14",
          5259 => x"3f",
          5260 => x"08",
          5261 => x"06",
          5262 => x"38",
          5263 => x"51",
          5264 => x"82",
          5265 => x"58",
          5266 => x"0c",
          5267 => x"33",
          5268 => x"80",
          5269 => x"ff",
          5270 => x"ff",
          5271 => x"55",
          5272 => x"81",
          5273 => x"38",
          5274 => x"06",
          5275 => x"fe",
          5276 => x"82",
          5277 => x"80",
          5278 => x"54",
          5279 => x"15",
          5280 => x"2e",
          5281 => x"13",
          5282 => x"72",
          5283 => x"38",
          5284 => x"ec",
          5285 => x"14",
          5286 => x"3f",
          5287 => x"08",
          5288 => x"ec",
          5289 => x"23",
          5290 => x"57",
          5291 => x"83",
          5292 => x"c7",
          5293 => x"ab",
          5294 => x"ec",
          5295 => x"ff",
          5296 => x"8d",
          5297 => x"14",
          5298 => x"3f",
          5299 => x"08",
          5300 => x"14",
          5301 => x"3f",
          5302 => x"08",
          5303 => x"06",
          5304 => x"79",
          5305 => x"98",
          5306 => x"22",
          5307 => x"84",
          5308 => x"5b",
          5309 => x"83",
          5310 => x"14",
          5311 => x"79",
          5312 => x"f8",
          5313 => x"85",
          5314 => x"82",
          5315 => x"80",
          5316 => x"38",
          5317 => x"08",
          5318 => x"ff",
          5319 => x"38",
          5320 => x"83",
          5321 => x"83",
          5322 => x"72",
          5323 => x"85",
          5324 => x"89",
          5325 => x"76",
          5326 => x"c4",
          5327 => x"70",
          5328 => x"7c",
          5329 => x"7a",
          5330 => x"17",
          5331 => x"ac",
          5332 => x"55",
          5333 => x"09",
          5334 => x"38",
          5335 => x"51",
          5336 => x"82",
          5337 => x"83",
          5338 => x"53",
          5339 => x"82",
          5340 => x"82",
          5341 => x"e0",
          5342 => x"fe",
          5343 => x"ec",
          5344 => x"0c",
          5345 => x"53",
          5346 => x"56",
          5347 => x"81",
          5348 => x"13",
          5349 => x"74",
          5350 => x"82",
          5351 => x"74",
          5352 => x"81",
          5353 => x"06",
          5354 => x"53",
          5355 => x"89",
          5356 => x"56",
          5357 => x"08",
          5358 => x"38",
          5359 => x"15",
          5360 => x"8c",
          5361 => x"80",
          5362 => x"34",
          5363 => x"09",
          5364 => x"92",
          5365 => x"14",
          5366 => x"3f",
          5367 => x"08",
          5368 => x"06",
          5369 => x"2e",
          5370 => x"80",
          5371 => x"1c",
          5372 => x"db",
          5373 => x"85",
          5374 => x"ea",
          5375 => x"ec",
          5376 => x"34",
          5377 => x"51",
          5378 => x"82",
          5379 => x"83",
          5380 => x"53",
          5381 => x"d5",
          5382 => x"06",
          5383 => x"b4",
          5384 => x"d6",
          5385 => x"ec",
          5386 => x"85",
          5387 => x"09",
          5388 => x"38",
          5389 => x"51",
          5390 => x"82",
          5391 => x"86",
          5392 => x"f2",
          5393 => x"06",
          5394 => x"9c",
          5395 => x"aa",
          5396 => x"ec",
          5397 => x"0c",
          5398 => x"51",
          5399 => x"82",
          5400 => x"8c",
          5401 => x"74",
          5402 => x"a0",
          5403 => x"53",
          5404 => x"a0",
          5405 => x"15",
          5406 => x"94",
          5407 => x"56",
          5408 => x"ec",
          5409 => x"0d",
          5410 => x"0d",
          5411 => x"55",
          5412 => x"b9",
          5413 => x"53",
          5414 => x"b1",
          5415 => x"52",
          5416 => x"a9",
          5417 => x"22",
          5418 => x"57",
          5419 => x"2e",
          5420 => x"99",
          5421 => x"33",
          5422 => x"3f",
          5423 => x"08",
          5424 => x"71",
          5425 => x"74",
          5426 => x"83",
          5427 => x"78",
          5428 => x"52",
          5429 => x"ec",
          5430 => x"0d",
          5431 => x"0d",
          5432 => x"33",
          5433 => x"3d",
          5434 => x"56",
          5435 => x"8b",
          5436 => x"82",
          5437 => x"24",
          5438 => x"85",
          5439 => x"2b",
          5440 => x"05",
          5441 => x"55",
          5442 => x"84",
          5443 => x"34",
          5444 => x"80",
          5445 => x"80",
          5446 => x"75",
          5447 => x"75",
          5448 => x"38",
          5449 => x"3d",
          5450 => x"05",
          5451 => x"3f",
          5452 => x"08",
          5453 => x"85",
          5454 => x"3d",
          5455 => x"3d",
          5456 => x"84",
          5457 => x"05",
          5458 => x"89",
          5459 => x"2e",
          5460 => x"77",
          5461 => x"54",
          5462 => x"05",
          5463 => x"84",
          5464 => x"f6",
          5465 => x"85",
          5466 => x"82",
          5467 => x"84",
          5468 => x"5c",
          5469 => x"3d",
          5470 => x"ed",
          5471 => x"85",
          5472 => x"82",
          5473 => x"92",
          5474 => x"d7",
          5475 => x"98",
          5476 => x"73",
          5477 => x"38",
          5478 => x"9c",
          5479 => x"80",
          5480 => x"38",
          5481 => x"95",
          5482 => x"2e",
          5483 => x"aa",
          5484 => x"ea",
          5485 => x"85",
          5486 => x"9e",
          5487 => x"05",
          5488 => x"54",
          5489 => x"38",
          5490 => x"70",
          5491 => x"54",
          5492 => x"8e",
          5493 => x"83",
          5494 => x"88",
          5495 => x"83",
          5496 => x"83",
          5497 => x"06",
          5498 => x"80",
          5499 => x"38",
          5500 => x"51",
          5501 => x"82",
          5502 => x"56",
          5503 => x"0a",
          5504 => x"05",
          5505 => x"3f",
          5506 => x"0b",
          5507 => x"80",
          5508 => x"7a",
          5509 => x"3f",
          5510 => x"9c",
          5511 => x"a3",
          5512 => x"81",
          5513 => x"34",
          5514 => x"80",
          5515 => x"b0",
          5516 => x"54",
          5517 => x"52",
          5518 => x"05",
          5519 => x"3f",
          5520 => x"08",
          5521 => x"ec",
          5522 => x"38",
          5523 => x"82",
          5524 => x"b2",
          5525 => x"84",
          5526 => x"06",
          5527 => x"73",
          5528 => x"38",
          5529 => x"af",
          5530 => x"2a",
          5531 => x"51",
          5532 => x"2e",
          5533 => x"81",
          5534 => x"80",
          5535 => x"87",
          5536 => x"39",
          5537 => x"51",
          5538 => x"82",
          5539 => x"7b",
          5540 => x"12",
          5541 => x"82",
          5542 => x"81",
          5543 => x"83",
          5544 => x"06",
          5545 => x"80",
          5546 => x"77",
          5547 => x"58",
          5548 => x"08",
          5549 => x"63",
          5550 => x"63",
          5551 => x"57",
          5552 => x"82",
          5553 => x"82",
          5554 => x"88",
          5555 => x"9c",
          5556 => x"d2",
          5557 => x"85",
          5558 => x"85",
          5559 => x"1b",
          5560 => x"0c",
          5561 => x"22",
          5562 => x"77",
          5563 => x"80",
          5564 => x"34",
          5565 => x"1a",
          5566 => x"94",
          5567 => x"85",
          5568 => x"06",
          5569 => x"80",
          5570 => x"38",
          5571 => x"08",
          5572 => x"86",
          5573 => x"ec",
          5574 => x"0c",
          5575 => x"70",
          5576 => x"52",
          5577 => x"39",
          5578 => x"51",
          5579 => x"82",
          5580 => x"57",
          5581 => x"08",
          5582 => x"38",
          5583 => x"85",
          5584 => x"2e",
          5585 => x"83",
          5586 => x"75",
          5587 => x"74",
          5588 => x"70",
          5589 => x"25",
          5590 => x"76",
          5591 => x"81",
          5592 => x"55",
          5593 => x"38",
          5594 => x"0c",
          5595 => x"75",
          5596 => x"54",
          5597 => x"a2",
          5598 => x"7a",
          5599 => x"3f",
          5600 => x"08",
          5601 => x"55",
          5602 => x"89",
          5603 => x"ec",
          5604 => x"1a",
          5605 => x"80",
          5606 => x"54",
          5607 => x"ec",
          5608 => x"0d",
          5609 => x"0d",
          5610 => x"64",
          5611 => x"59",
          5612 => x"90",
          5613 => x"52",
          5614 => x"cd",
          5615 => x"ec",
          5616 => x"85",
          5617 => x"38",
          5618 => x"55",
          5619 => x"86",
          5620 => x"82",
          5621 => x"19",
          5622 => x"55",
          5623 => x"80",
          5624 => x"38",
          5625 => x"0b",
          5626 => x"82",
          5627 => x"39",
          5628 => x"1a",
          5629 => x"82",
          5630 => x"19",
          5631 => x"08",
          5632 => x"7c",
          5633 => x"74",
          5634 => x"2e",
          5635 => x"94",
          5636 => x"83",
          5637 => x"56",
          5638 => x"38",
          5639 => x"22",
          5640 => x"89",
          5641 => x"55",
          5642 => x"75",
          5643 => x"19",
          5644 => x"39",
          5645 => x"52",
          5646 => x"ea",
          5647 => x"ec",
          5648 => x"75",
          5649 => x"38",
          5650 => x"ff",
          5651 => x"98",
          5652 => x"19",
          5653 => x"51",
          5654 => x"82",
          5655 => x"80",
          5656 => x"38",
          5657 => x"08",
          5658 => x"2a",
          5659 => x"80",
          5660 => x"38",
          5661 => x"8a",
          5662 => x"5c",
          5663 => x"27",
          5664 => x"7a",
          5665 => x"54",
          5666 => x"52",
          5667 => x"51",
          5668 => x"82",
          5669 => x"fe",
          5670 => x"83",
          5671 => x"56",
          5672 => x"9f",
          5673 => x"08",
          5674 => x"74",
          5675 => x"38",
          5676 => x"b4",
          5677 => x"16",
          5678 => x"89",
          5679 => x"51",
          5680 => x"77",
          5681 => x"b9",
          5682 => x"1a",
          5683 => x"08",
          5684 => x"84",
          5685 => x"57",
          5686 => x"27",
          5687 => x"56",
          5688 => x"52",
          5689 => x"97",
          5690 => x"ec",
          5691 => x"38",
          5692 => x"19",
          5693 => x"06",
          5694 => x"52",
          5695 => x"f2",
          5696 => x"31",
          5697 => x"7f",
          5698 => x"94",
          5699 => x"94",
          5700 => x"5c",
          5701 => x"80",
          5702 => x"85",
          5703 => x"3d",
          5704 => x"3d",
          5705 => x"65",
          5706 => x"5d",
          5707 => x"0c",
          5708 => x"05",
          5709 => x"f6",
          5710 => x"85",
          5711 => x"82",
          5712 => x"8a",
          5713 => x"33",
          5714 => x"2e",
          5715 => x"56",
          5716 => x"90",
          5717 => x"81",
          5718 => x"06",
          5719 => x"87",
          5720 => x"2e",
          5721 => x"95",
          5722 => x"91",
          5723 => x"56",
          5724 => x"81",
          5725 => x"34",
          5726 => x"8e",
          5727 => x"08",
          5728 => x"56",
          5729 => x"84",
          5730 => x"5c",
          5731 => x"82",
          5732 => x"18",
          5733 => x"ff",
          5734 => x"74",
          5735 => x"7e",
          5736 => x"ff",
          5737 => x"2a",
          5738 => x"7a",
          5739 => x"8c",
          5740 => x"08",
          5741 => x"38",
          5742 => x"39",
          5743 => x"52",
          5744 => x"be",
          5745 => x"ec",
          5746 => x"85",
          5747 => x"2e",
          5748 => x"74",
          5749 => x"91",
          5750 => x"2e",
          5751 => x"74",
          5752 => x"88",
          5753 => x"38",
          5754 => x"0c",
          5755 => x"15",
          5756 => x"08",
          5757 => x"06",
          5758 => x"51",
          5759 => x"82",
          5760 => x"fe",
          5761 => x"18",
          5762 => x"51",
          5763 => x"82",
          5764 => x"80",
          5765 => x"38",
          5766 => x"08",
          5767 => x"2a",
          5768 => x"80",
          5769 => x"38",
          5770 => x"8a",
          5771 => x"5b",
          5772 => x"27",
          5773 => x"7b",
          5774 => x"54",
          5775 => x"52",
          5776 => x"51",
          5777 => x"82",
          5778 => x"fe",
          5779 => x"b0",
          5780 => x"31",
          5781 => x"79",
          5782 => x"84",
          5783 => x"16",
          5784 => x"89",
          5785 => x"52",
          5786 => x"cc",
          5787 => x"55",
          5788 => x"16",
          5789 => x"2b",
          5790 => x"39",
          5791 => x"94",
          5792 => x"93",
          5793 => x"cd",
          5794 => x"85",
          5795 => x"e3",
          5796 => x"b0",
          5797 => x"76",
          5798 => x"94",
          5799 => x"ff",
          5800 => x"71",
          5801 => x"7b",
          5802 => x"38",
          5803 => x"18",
          5804 => x"51",
          5805 => x"82",
          5806 => x"fd",
          5807 => x"53",
          5808 => x"18",
          5809 => x"06",
          5810 => x"51",
          5811 => x"7e",
          5812 => x"83",
          5813 => x"76",
          5814 => x"17",
          5815 => x"1e",
          5816 => x"18",
          5817 => x"0c",
          5818 => x"58",
          5819 => x"74",
          5820 => x"38",
          5821 => x"8c",
          5822 => x"90",
          5823 => x"33",
          5824 => x"55",
          5825 => x"34",
          5826 => x"82",
          5827 => x"90",
          5828 => x"f8",
          5829 => x"8b",
          5830 => x"53",
          5831 => x"f2",
          5832 => x"85",
          5833 => x"82",
          5834 => x"80",
          5835 => x"16",
          5836 => x"2a",
          5837 => x"51",
          5838 => x"80",
          5839 => x"38",
          5840 => x"52",
          5841 => x"b7",
          5842 => x"ec",
          5843 => x"85",
          5844 => x"d4",
          5845 => x"08",
          5846 => x"a0",
          5847 => x"73",
          5848 => x"88",
          5849 => x"74",
          5850 => x"51",
          5851 => x"8c",
          5852 => x"9c",
          5853 => x"cb",
          5854 => x"b2",
          5855 => x"15",
          5856 => x"3f",
          5857 => x"15",
          5858 => x"3f",
          5859 => x"0b",
          5860 => x"78",
          5861 => x"3f",
          5862 => x"08",
          5863 => x"81",
          5864 => x"57",
          5865 => x"34",
          5866 => x"ec",
          5867 => x"0d",
          5868 => x"0d",
          5869 => x"54",
          5870 => x"82",
          5871 => x"53",
          5872 => x"08",
          5873 => x"3d",
          5874 => x"73",
          5875 => x"3f",
          5876 => x"08",
          5877 => x"ec",
          5878 => x"82",
          5879 => x"74",
          5880 => x"85",
          5881 => x"3d",
          5882 => x"3d",
          5883 => x"51",
          5884 => x"8b",
          5885 => x"82",
          5886 => x"24",
          5887 => x"85",
          5888 => x"9d",
          5889 => x"52",
          5890 => x"ec",
          5891 => x"0d",
          5892 => x"0d",
          5893 => x"3d",
          5894 => x"94",
          5895 => x"b8",
          5896 => x"ec",
          5897 => x"85",
          5898 => x"e0",
          5899 => x"63",
          5900 => x"d4",
          5901 => x"ec",
          5902 => x"ec",
          5903 => x"85",
          5904 => x"38",
          5905 => x"05",
          5906 => x"2b",
          5907 => x"80",
          5908 => x"76",
          5909 => x"0c",
          5910 => x"02",
          5911 => x"70",
          5912 => x"81",
          5913 => x"56",
          5914 => x"9e",
          5915 => x"53",
          5916 => x"db",
          5917 => x"85",
          5918 => x"15",
          5919 => x"82",
          5920 => x"84",
          5921 => x"06",
          5922 => x"55",
          5923 => x"ec",
          5924 => x"0d",
          5925 => x"0d",
          5926 => x"5b",
          5927 => x"80",
          5928 => x"ff",
          5929 => x"9f",
          5930 => x"ac",
          5931 => x"ec",
          5932 => x"85",
          5933 => x"fb",
          5934 => x"7a",
          5935 => x"08",
          5936 => x"64",
          5937 => x"2e",
          5938 => x"a0",
          5939 => x"70",
          5940 => x"c9",
          5941 => x"ec",
          5942 => x"85",
          5943 => x"d3",
          5944 => x"7b",
          5945 => x"3f",
          5946 => x"08",
          5947 => x"ec",
          5948 => x"38",
          5949 => x"51",
          5950 => x"82",
          5951 => x"45",
          5952 => x"51",
          5953 => x"82",
          5954 => x"57",
          5955 => x"08",
          5956 => x"80",
          5957 => x"da",
          5958 => x"85",
          5959 => x"82",
          5960 => x"a4",
          5961 => x"7b",
          5962 => x"3f",
          5963 => x"ec",
          5964 => x"38",
          5965 => x"51",
          5966 => x"82",
          5967 => x"57",
          5968 => x"08",
          5969 => x"38",
          5970 => x"09",
          5971 => x"38",
          5972 => x"df",
          5973 => x"db",
          5974 => x"ff",
          5975 => x"74",
          5976 => x"3f",
          5977 => x"78",
          5978 => x"33",
          5979 => x"56",
          5980 => x"91",
          5981 => x"05",
          5982 => x"81",
          5983 => x"56",
          5984 => x"f5",
          5985 => x"54",
          5986 => x"81",
          5987 => x"80",
          5988 => x"78",
          5989 => x"55",
          5990 => x"11",
          5991 => x"18",
          5992 => x"58",
          5993 => x"34",
          5994 => x"ff",
          5995 => x"55",
          5996 => x"34",
          5997 => x"77",
          5998 => x"81",
          5999 => x"ff",
          6000 => x"55",
          6001 => x"34",
          6002 => x"9d",
          6003 => x"82",
          6004 => x"a4",
          6005 => x"33",
          6006 => x"56",
          6007 => x"2e",
          6008 => x"16",
          6009 => x"33",
          6010 => x"73",
          6011 => x"16",
          6012 => x"26",
          6013 => x"55",
          6014 => x"91",
          6015 => x"54",
          6016 => x"70",
          6017 => x"34",
          6018 => x"ec",
          6019 => x"70",
          6020 => x"34",
          6021 => x"09",
          6022 => x"38",
          6023 => x"39",
          6024 => x"19",
          6025 => x"33",
          6026 => x"05",
          6027 => x"78",
          6028 => x"80",
          6029 => x"82",
          6030 => x"9e",
          6031 => x"f7",
          6032 => x"7d",
          6033 => x"05",
          6034 => x"57",
          6035 => x"3f",
          6036 => x"08",
          6037 => x"ec",
          6038 => x"38",
          6039 => x"53",
          6040 => x"38",
          6041 => x"54",
          6042 => x"92",
          6043 => x"33",
          6044 => x"70",
          6045 => x"54",
          6046 => x"38",
          6047 => x"15",
          6048 => x"70",
          6049 => x"58",
          6050 => x"82",
          6051 => x"8a",
          6052 => x"89",
          6053 => x"53",
          6054 => x"b9",
          6055 => x"ff",
          6056 => x"e0",
          6057 => x"85",
          6058 => x"15",
          6059 => x"53",
          6060 => x"e0",
          6061 => x"85",
          6062 => x"26",
          6063 => x"09",
          6064 => x"75",
          6065 => x"18",
          6066 => x"31",
          6067 => x"57",
          6068 => x"b1",
          6069 => x"08",
          6070 => x"38",
          6071 => x"51",
          6072 => x"82",
          6073 => x"54",
          6074 => x"08",
          6075 => x"9a",
          6076 => x"ec",
          6077 => x"81",
          6078 => x"85",
          6079 => x"16",
          6080 => x"16",
          6081 => x"2e",
          6082 => x"76",
          6083 => x"dc",
          6084 => x"31",
          6085 => x"18",
          6086 => x"90",
          6087 => x"81",
          6088 => x"06",
          6089 => x"56",
          6090 => x"9a",
          6091 => x"74",
          6092 => x"3f",
          6093 => x"08",
          6094 => x"ec",
          6095 => x"82",
          6096 => x"56",
          6097 => x"52",
          6098 => x"da",
          6099 => x"ec",
          6100 => x"ff",
          6101 => x"81",
          6102 => x"38",
          6103 => x"98",
          6104 => x"a6",
          6105 => x"16",
          6106 => x"39",
          6107 => x"16",
          6108 => x"75",
          6109 => x"53",
          6110 => x"aa",
          6111 => x"79",
          6112 => x"3f",
          6113 => x"08",
          6114 => x"0b",
          6115 => x"82",
          6116 => x"39",
          6117 => x"16",
          6118 => x"bb",
          6119 => x"2a",
          6120 => x"08",
          6121 => x"15",
          6122 => x"15",
          6123 => x"90",
          6124 => x"16",
          6125 => x"33",
          6126 => x"53",
          6127 => x"34",
          6128 => x"06",
          6129 => x"2e",
          6130 => x"9c",
          6131 => x"85",
          6132 => x"16",
          6133 => x"72",
          6134 => x"0c",
          6135 => x"04",
          6136 => x"79",
          6137 => x"75",
          6138 => x"8a",
          6139 => x"89",
          6140 => x"52",
          6141 => x"05",
          6142 => x"3f",
          6143 => x"08",
          6144 => x"ec",
          6145 => x"38",
          6146 => x"7a",
          6147 => x"d8",
          6148 => x"85",
          6149 => x"82",
          6150 => x"80",
          6151 => x"16",
          6152 => x"2b",
          6153 => x"74",
          6154 => x"86",
          6155 => x"84",
          6156 => x"06",
          6157 => x"73",
          6158 => x"38",
          6159 => x"52",
          6160 => x"b8",
          6161 => x"ec",
          6162 => x"0c",
          6163 => x"14",
          6164 => x"23",
          6165 => x"51",
          6166 => x"82",
          6167 => x"55",
          6168 => x"09",
          6169 => x"38",
          6170 => x"39",
          6171 => x"84",
          6172 => x"0c",
          6173 => x"82",
          6174 => x"89",
          6175 => x"fc",
          6176 => x"87",
          6177 => x"53",
          6178 => x"e7",
          6179 => x"85",
          6180 => x"38",
          6181 => x"08",
          6182 => x"3d",
          6183 => x"3d",
          6184 => x"89",
          6185 => x"54",
          6186 => x"54",
          6187 => x"82",
          6188 => x"53",
          6189 => x"08",
          6190 => x"74",
          6191 => x"85",
          6192 => x"73",
          6193 => x"3f",
          6194 => x"08",
          6195 => x"39",
          6196 => x"08",
          6197 => x"d3",
          6198 => x"85",
          6199 => x"82",
          6200 => x"84",
          6201 => x"06",
          6202 => x"53",
          6203 => x"85",
          6204 => x"38",
          6205 => x"51",
          6206 => x"72",
          6207 => x"ce",
          6208 => x"85",
          6209 => x"32",
          6210 => x"05",
          6211 => x"9f",
          6212 => x"85",
          6213 => x"51",
          6214 => x"72",
          6215 => x"0c",
          6216 => x"04",
          6217 => x"65",
          6218 => x"89",
          6219 => x"96",
          6220 => x"df",
          6221 => x"85",
          6222 => x"82",
          6223 => x"b2",
          6224 => x"75",
          6225 => x"3f",
          6226 => x"08",
          6227 => x"ec",
          6228 => x"02",
          6229 => x"33",
          6230 => x"55",
          6231 => x"25",
          6232 => x"55",
          6233 => x"80",
          6234 => x"76",
          6235 => x"d4",
          6236 => x"82",
          6237 => x"94",
          6238 => x"f0",
          6239 => x"65",
          6240 => x"53",
          6241 => x"05",
          6242 => x"51",
          6243 => x"82",
          6244 => x"5b",
          6245 => x"08",
          6246 => x"7c",
          6247 => x"08",
          6248 => x"fe",
          6249 => x"08",
          6250 => x"55",
          6251 => x"91",
          6252 => x"0c",
          6253 => x"81",
          6254 => x"39",
          6255 => x"ce",
          6256 => x"ec",
          6257 => x"55",
          6258 => x"2e",
          6259 => x"80",
          6260 => x"75",
          6261 => x"52",
          6262 => x"05",
          6263 => x"3f",
          6264 => x"08",
          6265 => x"38",
          6266 => x"08",
          6267 => x"38",
          6268 => x"08",
          6269 => x"70",
          6270 => x"08",
          6271 => x"7a",
          6272 => x"7f",
          6273 => x"54",
          6274 => x"77",
          6275 => x"80",
          6276 => x"15",
          6277 => x"ec",
          6278 => x"75",
          6279 => x"52",
          6280 => x"52",
          6281 => x"d7",
          6282 => x"ec",
          6283 => x"85",
          6284 => x"da",
          6285 => x"33",
          6286 => x"1a",
          6287 => x"54",
          6288 => x"09",
          6289 => x"38",
          6290 => x"ff",
          6291 => x"82",
          6292 => x"83",
          6293 => x"70",
          6294 => x"70",
          6295 => x"82",
          6296 => x"51",
          6297 => x"b4",
          6298 => x"bb",
          6299 => x"85",
          6300 => x"0a",
          6301 => x"81",
          6302 => x"25",
          6303 => x"59",
          6304 => x"75",
          6305 => x"7a",
          6306 => x"ff",
          6307 => x"7c",
          6308 => x"90",
          6309 => x"11",
          6310 => x"56",
          6311 => x"15",
          6312 => x"85",
          6313 => x"3d",
          6314 => x"3d",
          6315 => x"3d",
          6316 => x"70",
          6317 => x"d1",
          6318 => x"ec",
          6319 => x"85",
          6320 => x"a8",
          6321 => x"33",
          6322 => x"a0",
          6323 => x"33",
          6324 => x"70",
          6325 => x"55",
          6326 => x"73",
          6327 => x"8e",
          6328 => x"08",
          6329 => x"18",
          6330 => x"80",
          6331 => x"38",
          6332 => x"08",
          6333 => x"08",
          6334 => x"c3",
          6335 => x"85",
          6336 => x"88",
          6337 => x"80",
          6338 => x"17",
          6339 => x"51",
          6340 => x"3f",
          6341 => x"08",
          6342 => x"81",
          6343 => x"81",
          6344 => x"ec",
          6345 => x"09",
          6346 => x"38",
          6347 => x"39",
          6348 => x"77",
          6349 => x"ec",
          6350 => x"08",
          6351 => x"98",
          6352 => x"82",
          6353 => x"52",
          6354 => x"8a",
          6355 => x"ec",
          6356 => x"17",
          6357 => x"0c",
          6358 => x"80",
          6359 => x"73",
          6360 => x"75",
          6361 => x"38",
          6362 => x"34",
          6363 => x"82",
          6364 => x"89",
          6365 => x"e2",
          6366 => x"53",
          6367 => x"a4",
          6368 => x"3d",
          6369 => x"3f",
          6370 => x"08",
          6371 => x"ec",
          6372 => x"38",
          6373 => x"3d",
          6374 => x"3d",
          6375 => x"d1",
          6376 => x"85",
          6377 => x"82",
          6378 => x"81",
          6379 => x"80",
          6380 => x"70",
          6381 => x"81",
          6382 => x"56",
          6383 => x"81",
          6384 => x"98",
          6385 => x"74",
          6386 => x"38",
          6387 => x"05",
          6388 => x"06",
          6389 => x"55",
          6390 => x"38",
          6391 => x"51",
          6392 => x"82",
          6393 => x"74",
          6394 => x"81",
          6395 => x"56",
          6396 => x"80",
          6397 => x"54",
          6398 => x"08",
          6399 => x"2e",
          6400 => x"73",
          6401 => x"ec",
          6402 => x"52",
          6403 => x"52",
          6404 => x"3f",
          6405 => x"08",
          6406 => x"ec",
          6407 => x"38",
          6408 => x"08",
          6409 => x"cc",
          6410 => x"85",
          6411 => x"82",
          6412 => x"86",
          6413 => x"80",
          6414 => x"85",
          6415 => x"2e",
          6416 => x"85",
          6417 => x"c2",
          6418 => x"ce",
          6419 => x"85",
          6420 => x"85",
          6421 => x"81",
          6422 => x"85",
          6423 => x"80",
          6424 => x"55",
          6425 => x"94",
          6426 => x"2e",
          6427 => x"53",
          6428 => x"51",
          6429 => x"82",
          6430 => x"55",
          6431 => x"78",
          6432 => x"c2",
          6433 => x"ec",
          6434 => x"82",
          6435 => x"a0",
          6436 => x"e9",
          6437 => x"53",
          6438 => x"05",
          6439 => x"51",
          6440 => x"82",
          6441 => x"54",
          6442 => x"08",
          6443 => x"78",
          6444 => x"8e",
          6445 => x"58",
          6446 => x"82",
          6447 => x"54",
          6448 => x"08",
          6449 => x"54",
          6450 => x"82",
          6451 => x"84",
          6452 => x"06",
          6453 => x"02",
          6454 => x"33",
          6455 => x"81",
          6456 => x"86",
          6457 => x"f6",
          6458 => x"74",
          6459 => x"70",
          6460 => x"8e",
          6461 => x"ec",
          6462 => x"56",
          6463 => x"08",
          6464 => x"54",
          6465 => x"08",
          6466 => x"81",
          6467 => x"82",
          6468 => x"ec",
          6469 => x"09",
          6470 => x"38",
          6471 => x"b4",
          6472 => x"b0",
          6473 => x"ec",
          6474 => x"51",
          6475 => x"82",
          6476 => x"54",
          6477 => x"08",
          6478 => x"8b",
          6479 => x"b4",
          6480 => x"b6",
          6481 => x"54",
          6482 => x"15",
          6483 => x"90",
          6484 => x"34",
          6485 => x"0a",
          6486 => x"19",
          6487 => x"e3",
          6488 => x"78",
          6489 => x"51",
          6490 => x"a0",
          6491 => x"11",
          6492 => x"05",
          6493 => x"fa",
          6494 => x"ae",
          6495 => x"15",
          6496 => x"78",
          6497 => x"53",
          6498 => x"3f",
          6499 => x"0b",
          6500 => x"77",
          6501 => x"3f",
          6502 => x"08",
          6503 => x"ec",
          6504 => x"82",
          6505 => x"52",
          6506 => x"51",
          6507 => x"3f",
          6508 => x"52",
          6509 => x"fd",
          6510 => x"90",
          6511 => x"34",
          6512 => x"0b",
          6513 => x"78",
          6514 => x"fa",
          6515 => x"ec",
          6516 => x"39",
          6517 => x"52",
          6518 => x"bd",
          6519 => x"82",
          6520 => x"99",
          6521 => x"da",
          6522 => x"3d",
          6523 => x"d2",
          6524 => x"53",
          6525 => x"84",
          6526 => x"3d",
          6527 => x"3f",
          6528 => x"08",
          6529 => x"ec",
          6530 => x"38",
          6531 => x"3d",
          6532 => x"3d",
          6533 => x"cc",
          6534 => x"85",
          6535 => x"82",
          6536 => x"82",
          6537 => x"81",
          6538 => x"81",
          6539 => x"86",
          6540 => x"aa",
          6541 => x"a4",
          6542 => x"a8",
          6543 => x"05",
          6544 => x"ae",
          6545 => x"77",
          6546 => x"70",
          6547 => x"b4",
          6548 => x"3d",
          6549 => x"51",
          6550 => x"82",
          6551 => x"55",
          6552 => x"08",
          6553 => x"6f",
          6554 => x"06",
          6555 => x"a2",
          6556 => x"92",
          6557 => x"81",
          6558 => x"85",
          6559 => x"2e",
          6560 => x"81",
          6561 => x"51",
          6562 => x"82",
          6563 => x"55",
          6564 => x"08",
          6565 => x"68",
          6566 => x"a8",
          6567 => x"05",
          6568 => x"51",
          6569 => x"3f",
          6570 => x"33",
          6571 => x"8b",
          6572 => x"84",
          6573 => x"06",
          6574 => x"73",
          6575 => x"a0",
          6576 => x"8b",
          6577 => x"54",
          6578 => x"15",
          6579 => x"33",
          6580 => x"70",
          6581 => x"55",
          6582 => x"2e",
          6583 => x"6e",
          6584 => x"df",
          6585 => x"78",
          6586 => x"3f",
          6587 => x"08",
          6588 => x"ff",
          6589 => x"82",
          6590 => x"ec",
          6591 => x"80",
          6592 => x"85",
          6593 => x"78",
          6594 => x"f3",
          6595 => x"ec",
          6596 => x"d4",
          6597 => x"55",
          6598 => x"08",
          6599 => x"81",
          6600 => x"73",
          6601 => x"81",
          6602 => x"63",
          6603 => x"76",
          6604 => x"3f",
          6605 => x"0b",
          6606 => x"87",
          6607 => x"ec",
          6608 => x"77",
          6609 => x"3f",
          6610 => x"08",
          6611 => x"ec",
          6612 => x"78",
          6613 => x"ee",
          6614 => x"ec",
          6615 => x"82",
          6616 => x"a8",
          6617 => x"ed",
          6618 => x"80",
          6619 => x"02",
          6620 => x"df",
          6621 => x"57",
          6622 => x"3d",
          6623 => x"96",
          6624 => x"d4",
          6625 => x"ec",
          6626 => x"85",
          6627 => x"cf",
          6628 => x"65",
          6629 => x"d4",
          6630 => x"88",
          6631 => x"ec",
          6632 => x"85",
          6633 => x"38",
          6634 => x"05",
          6635 => x"06",
          6636 => x"73",
          6637 => x"a7",
          6638 => x"09",
          6639 => x"71",
          6640 => x"06",
          6641 => x"55",
          6642 => x"15",
          6643 => x"81",
          6644 => x"34",
          6645 => x"b3",
          6646 => x"85",
          6647 => x"74",
          6648 => x"0c",
          6649 => x"04",
          6650 => x"64",
          6651 => x"93",
          6652 => x"52",
          6653 => x"d1",
          6654 => x"85",
          6655 => x"82",
          6656 => x"80",
          6657 => x"58",
          6658 => x"3d",
          6659 => x"c8",
          6660 => x"85",
          6661 => x"82",
          6662 => x"b4",
          6663 => x"c7",
          6664 => x"a0",
          6665 => x"55",
          6666 => x"84",
          6667 => x"17",
          6668 => x"2b",
          6669 => x"96",
          6670 => x"b0",
          6671 => x"54",
          6672 => x"15",
          6673 => x"ff",
          6674 => x"82",
          6675 => x"55",
          6676 => x"ec",
          6677 => x"0d",
          6678 => x"0d",
          6679 => x"5a",
          6680 => x"3d",
          6681 => x"99",
          6682 => x"ec",
          6683 => x"ec",
          6684 => x"ec",
          6685 => x"05",
          6686 => x"ec",
          6687 => x"25",
          6688 => x"79",
          6689 => x"85",
          6690 => x"75",
          6691 => x"73",
          6692 => x"f9",
          6693 => x"80",
          6694 => x"8d",
          6695 => x"54",
          6696 => x"3f",
          6697 => x"08",
          6698 => x"ec",
          6699 => x"38",
          6700 => x"51",
          6701 => x"82",
          6702 => x"57",
          6703 => x"08",
          6704 => x"85",
          6705 => x"85",
          6706 => x"5b",
          6707 => x"18",
          6708 => x"18",
          6709 => x"74",
          6710 => x"81",
          6711 => x"78",
          6712 => x"8b",
          6713 => x"54",
          6714 => x"75",
          6715 => x"38",
          6716 => x"1b",
          6717 => x"55",
          6718 => x"2e",
          6719 => x"39",
          6720 => x"09",
          6721 => x"38",
          6722 => x"80",
          6723 => x"81",
          6724 => x"07",
          6725 => x"54",
          6726 => x"80",
          6727 => x"80",
          6728 => x"7b",
          6729 => x"53",
          6730 => x"d3",
          6731 => x"ec",
          6732 => x"85",
          6733 => x"38",
          6734 => x"55",
          6735 => x"56",
          6736 => x"8b",
          6737 => x"56",
          6738 => x"83",
          6739 => x"75",
          6740 => x"51",
          6741 => x"3f",
          6742 => x"08",
          6743 => x"82",
          6744 => x"98",
          6745 => x"e6",
          6746 => x"53",
          6747 => x"b8",
          6748 => x"3d",
          6749 => x"3f",
          6750 => x"08",
          6751 => x"08",
          6752 => x"85",
          6753 => x"98",
          6754 => x"a0",
          6755 => x"70",
          6756 => x"ae",
          6757 => x"6d",
          6758 => x"81",
          6759 => x"57",
          6760 => x"74",
          6761 => x"38",
          6762 => x"81",
          6763 => x"81",
          6764 => x"52",
          6765 => x"c9",
          6766 => x"ec",
          6767 => x"a5",
          6768 => x"33",
          6769 => x"54",
          6770 => x"3f",
          6771 => x"08",
          6772 => x"38",
          6773 => x"76",
          6774 => x"05",
          6775 => x"39",
          6776 => x"08",
          6777 => x"15",
          6778 => x"ff",
          6779 => x"73",
          6780 => x"38",
          6781 => x"83",
          6782 => x"56",
          6783 => x"75",
          6784 => x"81",
          6785 => x"33",
          6786 => x"2e",
          6787 => x"52",
          6788 => x"51",
          6789 => x"3f",
          6790 => x"08",
          6791 => x"ff",
          6792 => x"38",
          6793 => x"88",
          6794 => x"8a",
          6795 => x"38",
          6796 => x"ec",
          6797 => x"75",
          6798 => x"74",
          6799 => x"73",
          6800 => x"05",
          6801 => x"17",
          6802 => x"70",
          6803 => x"34",
          6804 => x"70",
          6805 => x"ff",
          6806 => x"55",
          6807 => x"26",
          6808 => x"8b",
          6809 => x"86",
          6810 => x"e5",
          6811 => x"38",
          6812 => x"99",
          6813 => x"05",
          6814 => x"70",
          6815 => x"73",
          6816 => x"81",
          6817 => x"ff",
          6818 => x"ed",
          6819 => x"80",
          6820 => x"91",
          6821 => x"55",
          6822 => x"3f",
          6823 => x"08",
          6824 => x"ec",
          6825 => x"38",
          6826 => x"51",
          6827 => x"3f",
          6828 => x"08",
          6829 => x"ec",
          6830 => x"76",
          6831 => x"67",
          6832 => x"34",
          6833 => x"82",
          6834 => x"84",
          6835 => x"06",
          6836 => x"80",
          6837 => x"2e",
          6838 => x"81",
          6839 => x"ff",
          6840 => x"82",
          6841 => x"54",
          6842 => x"08",
          6843 => x"53",
          6844 => x"08",
          6845 => x"ff",
          6846 => x"67",
          6847 => x"8b",
          6848 => x"53",
          6849 => x"51",
          6850 => x"3f",
          6851 => x"0b",
          6852 => x"79",
          6853 => x"ae",
          6854 => x"ec",
          6855 => x"55",
          6856 => x"ec",
          6857 => x"0d",
          6858 => x"0d",
          6859 => x"88",
          6860 => x"05",
          6861 => x"fc",
          6862 => x"54",
          6863 => x"d2",
          6864 => x"85",
          6865 => x"82",
          6866 => x"82",
          6867 => x"1a",
          6868 => x"82",
          6869 => x"80",
          6870 => x"8c",
          6871 => x"78",
          6872 => x"1a",
          6873 => x"2a",
          6874 => x"51",
          6875 => x"90",
          6876 => x"82",
          6877 => x"58",
          6878 => x"81",
          6879 => x"39",
          6880 => x"22",
          6881 => x"70",
          6882 => x"56",
          6883 => x"c6",
          6884 => x"14",
          6885 => x"09",
          6886 => x"72",
          6887 => x"82",
          6888 => x"05",
          6889 => x"7c",
          6890 => x"55",
          6891 => x"27",
          6892 => x"16",
          6893 => x"83",
          6894 => x"76",
          6895 => x"80",
          6896 => x"79",
          6897 => x"de",
          6898 => x"7f",
          6899 => x"14",
          6900 => x"83",
          6901 => x"82",
          6902 => x"81",
          6903 => x"38",
          6904 => x"08",
          6905 => x"93",
          6906 => x"ec",
          6907 => x"81",
          6908 => x"7b",
          6909 => x"06",
          6910 => x"39",
          6911 => x"56",
          6912 => x"09",
          6913 => x"b9",
          6914 => x"80",
          6915 => x"80",
          6916 => x"78",
          6917 => x"7a",
          6918 => x"38",
          6919 => x"73",
          6920 => x"81",
          6921 => x"ff",
          6922 => x"74",
          6923 => x"ff",
          6924 => x"82",
          6925 => x"58",
          6926 => x"08",
          6927 => x"74",
          6928 => x"16",
          6929 => x"73",
          6930 => x"39",
          6931 => x"7e",
          6932 => x"0c",
          6933 => x"2e",
          6934 => x"88",
          6935 => x"8c",
          6936 => x"1a",
          6937 => x"07",
          6938 => x"1b",
          6939 => x"08",
          6940 => x"16",
          6941 => x"75",
          6942 => x"38",
          6943 => x"90",
          6944 => x"15",
          6945 => x"54",
          6946 => x"34",
          6947 => x"82",
          6948 => x"90",
          6949 => x"e9",
          6950 => x"6d",
          6951 => x"80",
          6952 => x"9d",
          6953 => x"5c",
          6954 => x"3f",
          6955 => x"0b",
          6956 => x"08",
          6957 => x"38",
          6958 => x"08",
          6959 => x"9d",
          6960 => x"51",
          6961 => x"2e",
          6962 => x"75",
          6963 => x"ec",
          6964 => x"06",
          6965 => x"7e",
          6966 => x"8f",
          6967 => x"ec",
          6968 => x"06",
          6969 => x"56",
          6970 => x"74",
          6971 => x"76",
          6972 => x"81",
          6973 => x"8a",
          6974 => x"bd",
          6975 => x"fc",
          6976 => x"52",
          6977 => x"a4",
          6978 => x"85",
          6979 => x"38",
          6980 => x"80",
          6981 => x"74",
          6982 => x"26",
          6983 => x"15",
          6984 => x"74",
          6985 => x"38",
          6986 => x"80",
          6987 => x"84",
          6988 => x"92",
          6989 => x"80",
          6990 => x"38",
          6991 => x"06",
          6992 => x"2e",
          6993 => x"56",
          6994 => x"78",
          6995 => x"89",
          6996 => x"2b",
          6997 => x"43",
          6998 => x"38",
          6999 => x"09",
          7000 => x"80",
          7001 => x"51",
          7002 => x"74",
          7003 => x"99",
          7004 => x"53",
          7005 => x"51",
          7006 => x"3f",
          7007 => x"85",
          7008 => x"b5",
          7009 => x"2a",
          7010 => x"82",
          7011 => x"43",
          7012 => x"83",
          7013 => x"66",
          7014 => x"60",
          7015 => x"99",
          7016 => x"31",
          7017 => x"80",
          7018 => x"8a",
          7019 => x"56",
          7020 => x"26",
          7021 => x"77",
          7022 => x"81",
          7023 => x"74",
          7024 => x"38",
          7025 => x"55",
          7026 => x"83",
          7027 => x"81",
          7028 => x"80",
          7029 => x"38",
          7030 => x"55",
          7031 => x"5e",
          7032 => x"89",
          7033 => x"5a",
          7034 => x"09",
          7035 => x"e0",
          7036 => x"38",
          7037 => x"57",
          7038 => x"80",
          7039 => x"5a",
          7040 => x"9d",
          7041 => x"26",
          7042 => x"80",
          7043 => x"10",
          7044 => x"22",
          7045 => x"74",
          7046 => x"38",
          7047 => x"ee",
          7048 => x"66",
          7049 => x"e4",
          7050 => x"ec",
          7051 => x"84",
          7052 => x"2a",
          7053 => x"5c",
          7054 => x"85",
          7055 => x"80",
          7056 => x"44",
          7057 => x"0a",
          7058 => x"f2",
          7059 => x"39",
          7060 => x"66",
          7061 => x"81",
          7062 => x"c8",
          7063 => x"74",
          7064 => x"38",
          7065 => x"98",
          7066 => x"c8",
          7067 => x"82",
          7068 => x"57",
          7069 => x"80",
          7070 => x"76",
          7071 => x"38",
          7072 => x"51",
          7073 => x"3f",
          7074 => x"08",
          7075 => x"08",
          7076 => x"57",
          7077 => x"08",
          7078 => x"98",
          7079 => x"82",
          7080 => x"71",
          7081 => x"ec",
          7082 => x"70",
          7083 => x"05",
          7084 => x"5e",
          7085 => x"89",
          7086 => x"5c",
          7087 => x"1c",
          7088 => x"05",
          7089 => x"ff",
          7090 => x"81",
          7091 => x"06",
          7092 => x"52",
          7093 => x"40",
          7094 => x"09",
          7095 => x"38",
          7096 => x"18",
          7097 => x"39",
          7098 => x"79",
          7099 => x"19",
          7100 => x"58",
          7101 => x"76",
          7102 => x"38",
          7103 => x"7d",
          7104 => x"70",
          7105 => x"55",
          7106 => x"3f",
          7107 => x"08",
          7108 => x"2e",
          7109 => x"9b",
          7110 => x"ec",
          7111 => x"f5",
          7112 => x"38",
          7113 => x"38",
          7114 => x"59",
          7115 => x"38",
          7116 => x"7d",
          7117 => x"81",
          7118 => x"38",
          7119 => x"0b",
          7120 => x"08",
          7121 => x"78",
          7122 => x"1a",
          7123 => x"c0",
          7124 => x"74",
          7125 => x"39",
          7126 => x"55",
          7127 => x"8f",
          7128 => x"fd",
          7129 => x"85",
          7130 => x"f5",
          7131 => x"78",
          7132 => x"79",
          7133 => x"80",
          7134 => x"ea",
          7135 => x"39",
          7136 => x"81",
          7137 => x"06",
          7138 => x"55",
          7139 => x"27",
          7140 => x"81",
          7141 => x"56",
          7142 => x"38",
          7143 => x"80",
          7144 => x"ff",
          7145 => x"8b",
          7146 => x"f0",
          7147 => x"ff",
          7148 => x"84",
          7149 => x"1b",
          7150 => x"e9",
          7151 => x"1c",
          7152 => x"ff",
          7153 => x"8e",
          7154 => x"a0",
          7155 => x"0b",
          7156 => x"7d",
          7157 => x"09",
          7158 => x"96",
          7159 => x"06",
          7160 => x"91",
          7161 => x"a0",
          7162 => x"55",
          7163 => x"ff",
          7164 => x"74",
          7165 => x"06",
          7166 => x"51",
          7167 => x"3f",
          7168 => x"52",
          7169 => x"ff",
          7170 => x"f8",
          7171 => x"34",
          7172 => x"1b",
          7173 => x"8d",
          7174 => x"52",
          7175 => x"ff",
          7176 => x"60",
          7177 => x"51",
          7178 => x"3f",
          7179 => x"09",
          7180 => x"cb",
          7181 => x"b2",
          7182 => x"c3",
          7183 => x"a0",
          7184 => x"52",
          7185 => x"ff",
          7186 => x"82",
          7187 => x"51",
          7188 => x"3f",
          7189 => x"1b",
          7190 => x"c9",
          7191 => x"b2",
          7192 => x"9f",
          7193 => x"80",
          7194 => x"1c",
          7195 => x"80",
          7196 => x"93",
          7197 => x"fc",
          7198 => x"1b",
          7199 => x"82",
          7200 => x"52",
          7201 => x"ff",
          7202 => x"7c",
          7203 => x"06",
          7204 => x"51",
          7205 => x"3f",
          7206 => x"a4",
          7207 => x"0b",
          7208 => x"93",
          7209 => x"90",
          7210 => x"51",
          7211 => x"3f",
          7212 => x"52",
          7213 => x"70",
          7214 => x"9e",
          7215 => x"54",
          7216 => x"52",
          7217 => x"9b",
          7218 => x"56",
          7219 => x"08",
          7220 => x"7d",
          7221 => x"81",
          7222 => x"38",
          7223 => x"86",
          7224 => x"52",
          7225 => x"9a",
          7226 => x"80",
          7227 => x"7a",
          7228 => x"a1",
          7229 => x"85",
          7230 => x"7a",
          7231 => x"c3",
          7232 => x"85",
          7233 => x"83",
          7234 => x"ff",
          7235 => x"ff",
          7236 => x"e8",
          7237 => x"9e",
          7238 => x"52",
          7239 => x"51",
          7240 => x"3f",
          7241 => x"52",
          7242 => x"9d",
          7243 => x"54",
          7244 => x"53",
          7245 => x"51",
          7246 => x"3f",
          7247 => x"16",
          7248 => x"7e",
          7249 => x"8c",
          7250 => x"80",
          7251 => x"ff",
          7252 => x"7f",
          7253 => x"7d",
          7254 => x"81",
          7255 => x"f8",
          7256 => x"ff",
          7257 => x"ff",
          7258 => x"51",
          7259 => x"3f",
          7260 => x"88",
          7261 => x"39",
          7262 => x"f8",
          7263 => x"2e",
          7264 => x"55",
          7265 => x"51",
          7266 => x"3f",
          7267 => x"57",
          7268 => x"83",
          7269 => x"76",
          7270 => x"7a",
          7271 => x"ff",
          7272 => x"82",
          7273 => x"82",
          7274 => x"80",
          7275 => x"ec",
          7276 => x"51",
          7277 => x"3f",
          7278 => x"78",
          7279 => x"74",
          7280 => x"18",
          7281 => x"2e",
          7282 => x"79",
          7283 => x"2e",
          7284 => x"55",
          7285 => x"62",
          7286 => x"74",
          7287 => x"75",
          7288 => x"7e",
          7289 => x"ec",
          7290 => x"ec",
          7291 => x"38",
          7292 => x"78",
          7293 => x"74",
          7294 => x"56",
          7295 => x"93",
          7296 => x"66",
          7297 => x"26",
          7298 => x"56",
          7299 => x"83",
          7300 => x"64",
          7301 => x"77",
          7302 => x"84",
          7303 => x"52",
          7304 => x"9c",
          7305 => x"d4",
          7306 => x"51",
          7307 => x"3f",
          7308 => x"55",
          7309 => x"81",
          7310 => x"34",
          7311 => x"16",
          7312 => x"16",
          7313 => x"16",
          7314 => x"05",
          7315 => x"c1",
          7316 => x"fe",
          7317 => x"fe",
          7318 => x"34",
          7319 => x"08",
          7320 => x"07",
          7321 => x"16",
          7322 => x"ec",
          7323 => x"34",
          7324 => x"c6",
          7325 => x"9b",
          7326 => x"52",
          7327 => x"51",
          7328 => x"3f",
          7329 => x"53",
          7330 => x"51",
          7331 => x"3f",
          7332 => x"85",
          7333 => x"38",
          7334 => x"52",
          7335 => x"99",
          7336 => x"56",
          7337 => x"08",
          7338 => x"39",
          7339 => x"39",
          7340 => x"39",
          7341 => x"08",
          7342 => x"85",
          7343 => x"3d",
          7344 => x"3d",
          7345 => x"5b",
          7346 => x"60",
          7347 => x"57",
          7348 => x"25",
          7349 => x"3d",
          7350 => x"55",
          7351 => x"15",
          7352 => x"c9",
          7353 => x"81",
          7354 => x"06",
          7355 => x"3d",
          7356 => x"8d",
          7357 => x"74",
          7358 => x"05",
          7359 => x"17",
          7360 => x"2e",
          7361 => x"c9",
          7362 => x"34",
          7363 => x"83",
          7364 => x"74",
          7365 => x"0c",
          7366 => x"04",
          7367 => x"7b",
          7368 => x"b3",
          7369 => x"57",
          7370 => x"09",
          7371 => x"38",
          7372 => x"51",
          7373 => x"17",
          7374 => x"76",
          7375 => x"38",
          7376 => x"77",
          7377 => x"56",
          7378 => x"34",
          7379 => x"bb",
          7380 => x"38",
          7381 => x"05",
          7382 => x"8c",
          7383 => x"08",
          7384 => x"3f",
          7385 => x"70",
          7386 => x"70",
          7387 => x"2a",
          7388 => x"05",
          7389 => x"56",
          7390 => x"0c",
          7391 => x"18",
          7392 => x"0d",
          7393 => x"0d",
          7394 => x"08",
          7395 => x"75",
          7396 => x"89",
          7397 => x"54",
          7398 => x"16",
          7399 => x"51",
          7400 => x"82",
          7401 => x"91",
          7402 => x"08",
          7403 => x"81",
          7404 => x"88",
          7405 => x"83",
          7406 => x"74",
          7407 => x"0c",
          7408 => x"04",
          7409 => x"75",
          7410 => x"53",
          7411 => x"51",
          7412 => x"3f",
          7413 => x"85",
          7414 => x"ea",
          7415 => x"80",
          7416 => x"6a",
          7417 => x"70",
          7418 => x"d8",
          7419 => x"72",
          7420 => x"3f",
          7421 => x"8d",
          7422 => x"0d",
          7423 => x"ff",
          7424 => x"00",
          7425 => x"ff",
          7426 => x"ff",
          7427 => x"00",
          7428 => x"00",
          7429 => x"00",
          7430 => x"00",
          7431 => x"00",
          7432 => x"00",
          7433 => x"00",
          7434 => x"00",
          7435 => x"00",
          7436 => x"00",
          7437 => x"00",
          7438 => x"00",
          7439 => x"00",
          7440 => x"00",
          7441 => x"00",
          7442 => x"00",
          7443 => x"00",
          7444 => x"00",
          7445 => x"00",
          7446 => x"00",
          7447 => x"00",
          7448 => x"00",
          7449 => x"00",
          7450 => x"00",
          7451 => x"00",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"00",
          7462 => x"00",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"00",
          7467 => x"00",
          7468 => x"00",
          7469 => x"00",
          7470 => x"00",
          7471 => x"00",
          7472 => x"00",
          7473 => x"00",
          7474 => x"69",
          7475 => x"00",
          7476 => x"69",
          7477 => x"6c",
          7478 => x"69",
          7479 => x"00",
          7480 => x"6c",
          7481 => x"00",
          7482 => x"65",
          7483 => x"00",
          7484 => x"63",
          7485 => x"72",
          7486 => x"63",
          7487 => x"00",
          7488 => x"64",
          7489 => x"00",
          7490 => x"64",
          7491 => x"00",
          7492 => x"65",
          7493 => x"65",
          7494 => x"65",
          7495 => x"69",
          7496 => x"69",
          7497 => x"66",
          7498 => x"66",
          7499 => x"61",
          7500 => x"00",
          7501 => x"6d",
          7502 => x"65",
          7503 => x"72",
          7504 => x"65",
          7505 => x"00",
          7506 => x"6e",
          7507 => x"00",
          7508 => x"65",
          7509 => x"00",
          7510 => x"62",
          7511 => x"63",
          7512 => x"62",
          7513 => x"63",
          7514 => x"69",
          7515 => x"00",
          7516 => x"64",
          7517 => x"69",
          7518 => x"45",
          7519 => x"72",
          7520 => x"6e",
          7521 => x"6e",
          7522 => x"65",
          7523 => x"72",
          7524 => x"00",
          7525 => x"69",
          7526 => x"6e",
          7527 => x"72",
          7528 => x"79",
          7529 => x"00",
          7530 => x"6f",
          7531 => x"6c",
          7532 => x"6f",
          7533 => x"2e",
          7534 => x"6f",
          7535 => x"74",
          7536 => x"6f",
          7537 => x"2e",
          7538 => x"6e",
          7539 => x"69",
          7540 => x"69",
          7541 => x"61",
          7542 => x"0a",
          7543 => x"63",
          7544 => x"73",
          7545 => x"6e",
          7546 => x"2e",
          7547 => x"69",
          7548 => x"61",
          7549 => x"61",
          7550 => x"65",
          7551 => x"74",
          7552 => x"00",
          7553 => x"69",
          7554 => x"68",
          7555 => x"6c",
          7556 => x"6e",
          7557 => x"69",
          7558 => x"00",
          7559 => x"44",
          7560 => x"20",
          7561 => x"74",
          7562 => x"72",
          7563 => x"63",
          7564 => x"2e",
          7565 => x"72",
          7566 => x"20",
          7567 => x"62",
          7568 => x"69",
          7569 => x"6e",
          7570 => x"69",
          7571 => x"00",
          7572 => x"69",
          7573 => x"6e",
          7574 => x"65",
          7575 => x"6c",
          7576 => x"0a",
          7577 => x"6f",
          7578 => x"6d",
          7579 => x"69",
          7580 => x"20",
          7581 => x"65",
          7582 => x"74",
          7583 => x"66",
          7584 => x"64",
          7585 => x"20",
          7586 => x"6b",
          7587 => x"00",
          7588 => x"6f",
          7589 => x"74",
          7590 => x"6f",
          7591 => x"64",
          7592 => x"00",
          7593 => x"69",
          7594 => x"75",
          7595 => x"6f",
          7596 => x"61",
          7597 => x"6e",
          7598 => x"6e",
          7599 => x"6c",
          7600 => x"0a",
          7601 => x"69",
          7602 => x"69",
          7603 => x"6f",
          7604 => x"64",
          7605 => x"00",
          7606 => x"6e",
          7607 => x"66",
          7608 => x"65",
          7609 => x"6d",
          7610 => x"72",
          7611 => x"00",
          7612 => x"6f",
          7613 => x"61",
          7614 => x"6f",
          7615 => x"20",
          7616 => x"65",
          7617 => x"00",
          7618 => x"61",
          7619 => x"65",
          7620 => x"73",
          7621 => x"63",
          7622 => x"65",
          7623 => x"0a",
          7624 => x"75",
          7625 => x"73",
          7626 => x"00",
          7627 => x"6e",
          7628 => x"77",
          7629 => x"72",
          7630 => x"2e",
          7631 => x"25",
          7632 => x"62",
          7633 => x"73",
          7634 => x"20",
          7635 => x"25",
          7636 => x"62",
          7637 => x"73",
          7638 => x"63",
          7639 => x"00",
          7640 => x"65",
          7641 => x"00",
          7642 => x"30",
          7643 => x"00",
          7644 => x"20",
          7645 => x"30",
          7646 => x"00",
          7647 => x"20",
          7648 => x"20",
          7649 => x"00",
          7650 => x"30",
          7651 => x"00",
          7652 => x"20",
          7653 => x"7c",
          7654 => x"0d",
          7655 => x"4f",
          7656 => x"2a",
          7657 => x"73",
          7658 => x"00",
          7659 => x"32",
          7660 => x"2f",
          7661 => x"30",
          7662 => x"31",
          7663 => x"00",
          7664 => x"5a",
          7665 => x"20",
          7666 => x"20",
          7667 => x"78",
          7668 => x"73",
          7669 => x"20",
          7670 => x"0a",
          7671 => x"50",
          7672 => x"6e",
          7673 => x"72",
          7674 => x"20",
          7675 => x"64",
          7676 => x"0a",
          7677 => x"69",
          7678 => x"20",
          7679 => x"65",
          7680 => x"70",
          7681 => x"00",
          7682 => x"53",
          7683 => x"6e",
          7684 => x"72",
          7685 => x"0a",
          7686 => x"4f",
          7687 => x"20",
          7688 => x"69",
          7689 => x"72",
          7690 => x"74",
          7691 => x"4f",
          7692 => x"20",
          7693 => x"69",
          7694 => x"72",
          7695 => x"74",
          7696 => x"41",
          7697 => x"20",
          7698 => x"69",
          7699 => x"72",
          7700 => x"74",
          7701 => x"41",
          7702 => x"20",
          7703 => x"69",
          7704 => x"72",
          7705 => x"74",
          7706 => x"41",
          7707 => x"20",
          7708 => x"69",
          7709 => x"72",
          7710 => x"74",
          7711 => x"41",
          7712 => x"20",
          7713 => x"69",
          7714 => x"72",
          7715 => x"74",
          7716 => x"65",
          7717 => x"6e",
          7718 => x"70",
          7719 => x"6d",
          7720 => x"2e",
          7721 => x"00",
          7722 => x"6e",
          7723 => x"69",
          7724 => x"74",
          7725 => x"72",
          7726 => x"0a",
          7727 => x"75",
          7728 => x"78",
          7729 => x"62",
          7730 => x"00",
          7731 => x"4f",
          7732 => x"73",
          7733 => x"3a",
          7734 => x"61",
          7735 => x"64",
          7736 => x"20",
          7737 => x"74",
          7738 => x"69",
          7739 => x"73",
          7740 => x"61",
          7741 => x"30",
          7742 => x"6c",
          7743 => x"65",
          7744 => x"69",
          7745 => x"61",
          7746 => x"6c",
          7747 => x"0a",
          7748 => x"20",
          7749 => x"6c",
          7750 => x"69",
          7751 => x"2e",
          7752 => x"00",
          7753 => x"6f",
          7754 => x"6e",
          7755 => x"2e",
          7756 => x"6f",
          7757 => x"72",
          7758 => x"2e",
          7759 => x"00",
          7760 => x"30",
          7761 => x"28",
          7762 => x"78",
          7763 => x"25",
          7764 => x"78",
          7765 => x"38",
          7766 => x"00",
          7767 => x"75",
          7768 => x"4d",
          7769 => x"72",
          7770 => x"00",
          7771 => x"43",
          7772 => x"6c",
          7773 => x"2e",
          7774 => x"30",
          7775 => x"25",
          7776 => x"2d",
          7777 => x"3f",
          7778 => x"00",
          7779 => x"30",
          7780 => x"25",
          7781 => x"2d",
          7782 => x"30",
          7783 => x"25",
          7784 => x"2d",
          7785 => x"78",
          7786 => x"74",
          7787 => x"20",
          7788 => x"65",
          7789 => x"25",
          7790 => x"20",
          7791 => x"0a",
          7792 => x"61",
          7793 => x"6e",
          7794 => x"6f",
          7795 => x"40",
          7796 => x"38",
          7797 => x"2e",
          7798 => x"00",
          7799 => x"61",
          7800 => x"72",
          7801 => x"72",
          7802 => x"20",
          7803 => x"65",
          7804 => x"64",
          7805 => x"00",
          7806 => x"65",
          7807 => x"72",
          7808 => x"67",
          7809 => x"70",
          7810 => x"61",
          7811 => x"6e",
          7812 => x"0a",
          7813 => x"6f",
          7814 => x"72",
          7815 => x"6f",
          7816 => x"67",
          7817 => x"0a",
          7818 => x"50",
          7819 => x"69",
          7820 => x"64",
          7821 => x"73",
          7822 => x"2e",
          7823 => x"00",
          7824 => x"64",
          7825 => x"73",
          7826 => x"00",
          7827 => x"64",
          7828 => x"73",
          7829 => x"61",
          7830 => x"6f",
          7831 => x"6e",
          7832 => x"00",
          7833 => x"75",
          7834 => x"6e",
          7835 => x"2e",
          7836 => x"6e",
          7837 => x"69",
          7838 => x"69",
          7839 => x"72",
          7840 => x"74",
          7841 => x"2e",
          7842 => x"64",
          7843 => x"2f",
          7844 => x"25",
          7845 => x"64",
          7846 => x"2e",
          7847 => x"64",
          7848 => x"6f",
          7849 => x"6f",
          7850 => x"67",
          7851 => x"74",
          7852 => x"00",
          7853 => x"28",
          7854 => x"6d",
          7855 => x"43",
          7856 => x"6e",
          7857 => x"29",
          7858 => x"0a",
          7859 => x"69",
          7860 => x"20",
          7861 => x"6c",
          7862 => x"6e",
          7863 => x"3a",
          7864 => x"20",
          7865 => x"42",
          7866 => x"52",
          7867 => x"20",
          7868 => x"38",
          7869 => x"30",
          7870 => x"2e",
          7871 => x"20",
          7872 => x"44",
          7873 => x"20",
          7874 => x"20",
          7875 => x"38",
          7876 => x"30",
          7877 => x"2e",
          7878 => x"20",
          7879 => x"4e",
          7880 => x"42",
          7881 => x"20",
          7882 => x"38",
          7883 => x"30",
          7884 => x"2e",
          7885 => x"20",
          7886 => x"52",
          7887 => x"20",
          7888 => x"20",
          7889 => x"38",
          7890 => x"30",
          7891 => x"2e",
          7892 => x"20",
          7893 => x"41",
          7894 => x"20",
          7895 => x"20",
          7896 => x"38",
          7897 => x"30",
          7898 => x"2e",
          7899 => x"20",
          7900 => x"44",
          7901 => x"52",
          7902 => x"20",
          7903 => x"76",
          7904 => x"73",
          7905 => x"30",
          7906 => x"2e",
          7907 => x"20",
          7908 => x"49",
          7909 => x"31",
          7910 => x"20",
          7911 => x"6d",
          7912 => x"20",
          7913 => x"30",
          7914 => x"2e",
          7915 => x"20",
          7916 => x"4e",
          7917 => x"43",
          7918 => x"20",
          7919 => x"61",
          7920 => x"6c",
          7921 => x"30",
          7922 => x"2e",
          7923 => x"20",
          7924 => x"49",
          7925 => x"4f",
          7926 => x"42",
          7927 => x"00",
          7928 => x"20",
          7929 => x"42",
          7930 => x"43",
          7931 => x"20",
          7932 => x"4f",
          7933 => x"0a",
          7934 => x"20",
          7935 => x"53",
          7936 => x"00",
          7937 => x"20",
          7938 => x"50",
          7939 => x"00",
          7940 => x"64",
          7941 => x"73",
          7942 => x"3a",
          7943 => x"20",
          7944 => x"50",
          7945 => x"65",
          7946 => x"20",
          7947 => x"74",
          7948 => x"41",
          7949 => x"65",
          7950 => x"3d",
          7951 => x"38",
          7952 => x"00",
          7953 => x"20",
          7954 => x"50",
          7955 => x"65",
          7956 => x"79",
          7957 => x"61",
          7958 => x"41",
          7959 => x"65",
          7960 => x"3d",
          7961 => x"38",
          7962 => x"00",
          7963 => x"20",
          7964 => x"74",
          7965 => x"20",
          7966 => x"72",
          7967 => x"64",
          7968 => x"73",
          7969 => x"20",
          7970 => x"3d",
          7971 => x"38",
          7972 => x"00",
          7973 => x"69",
          7974 => x"0a",
          7975 => x"20",
          7976 => x"50",
          7977 => x"64",
          7978 => x"20",
          7979 => x"20",
          7980 => x"20",
          7981 => x"20",
          7982 => x"3d",
          7983 => x"34",
          7984 => x"00",
          7985 => x"20",
          7986 => x"79",
          7987 => x"6d",
          7988 => x"6f",
          7989 => x"46",
          7990 => x"20",
          7991 => x"20",
          7992 => x"3d",
          7993 => x"2e",
          7994 => x"64",
          7995 => x"0a",
          7996 => x"20",
          7997 => x"44",
          7998 => x"20",
          7999 => x"63",
          8000 => x"72",
          8001 => x"20",
          8002 => x"20",
          8003 => x"3d",
          8004 => x"2e",
          8005 => x"64",
          8006 => x"0a",
          8007 => x"20",
          8008 => x"69",
          8009 => x"6f",
          8010 => x"53",
          8011 => x"4d",
          8012 => x"6f",
          8013 => x"46",
          8014 => x"3d",
          8015 => x"2e",
          8016 => x"64",
          8017 => x"0a",
          8018 => x"6d",
          8019 => x"00",
          8020 => x"65",
          8021 => x"6d",
          8022 => x"6c",
          8023 => x"00",
          8024 => x"56",
          8025 => x"56",
          8026 => x"6e",
          8027 => x"6e",
          8028 => x"77",
          8029 => x"00",
          8030 => x"00",
          8031 => x"00",
          8032 => x"00",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"5b",
          8096 => x"5b",
          8097 => x"5b",
          8098 => x"5b",
          8099 => x"5b",
          8100 => x"5b",
          8101 => x"5b",
          8102 => x"30",
          8103 => x"5b",
          8104 => x"5b",
          8105 => x"5b",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"69",
          8118 => x"72",
          8119 => x"69",
          8120 => x"00",
          8121 => x"00",
          8122 => x"30",
          8123 => x"20",
          8124 => x"00",
          8125 => x"61",
          8126 => x"64",
          8127 => x"20",
          8128 => x"65",
          8129 => x"68",
          8130 => x"69",
          8131 => x"72",
          8132 => x"69",
          8133 => x"74",
          8134 => x"4f",
          8135 => x"00",
          8136 => x"61",
          8137 => x"74",
          8138 => x"65",
          8139 => x"72",
          8140 => x"65",
          8141 => x"73",
          8142 => x"79",
          8143 => x"6c",
          8144 => x"64",
          8145 => x"62",
          8146 => x"67",
          8147 => x"00",
          8148 => x"44",
          8149 => x"2a",
          8150 => x"3b",
          8151 => x"3f",
          8152 => x"7f",
          8153 => x"41",
          8154 => x"41",
          8155 => x"00",
          8156 => x"fe",
          8157 => x"44",
          8158 => x"2e",
          8159 => x"4f",
          8160 => x"4d",
          8161 => x"20",
          8162 => x"54",
          8163 => x"20",
          8164 => x"4f",
          8165 => x"4d",
          8166 => x"20",
          8167 => x"54",
          8168 => x"20",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"9a",
          8174 => x"41",
          8175 => x"45",
          8176 => x"49",
          8177 => x"92",
          8178 => x"4f",
          8179 => x"99",
          8180 => x"9d",
          8181 => x"49",
          8182 => x"a5",
          8183 => x"a9",
          8184 => x"ad",
          8185 => x"b1",
          8186 => x"b5",
          8187 => x"b9",
          8188 => x"bd",
          8189 => x"c1",
          8190 => x"c5",
          8191 => x"c9",
          8192 => x"cd",
          8193 => x"d1",
          8194 => x"d5",
          8195 => x"d9",
          8196 => x"dd",
          8197 => x"e1",
          8198 => x"e5",
          8199 => x"e9",
          8200 => x"ed",
          8201 => x"f1",
          8202 => x"f5",
          8203 => x"f9",
          8204 => x"fd",
          8205 => x"2e",
          8206 => x"5b",
          8207 => x"22",
          8208 => x"3e",
          8209 => x"00",
          8210 => x"01",
          8211 => x"10",
          8212 => x"00",
          8213 => x"00",
          8214 => x"01",
          8215 => x"04",
          8216 => x"10",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"02",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"04",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"14",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"2b",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"30",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"3c",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"3d",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"3f",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"40",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"41",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"42",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"43",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"50",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"51",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"54",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"55",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"79",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"78",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"82",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"83",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"85",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"87",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"8c",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"8d",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"8e",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"8f",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"01",
          8329 => x"00",
          8330 => x"01",
          8331 => x"81",
          8332 => x"00",
          8333 => x"7f",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"f5",
          8339 => x"f5",
          8340 => x"f5",
          8341 => x"00",
          8342 => x"01",
          8343 => x"01",
          8344 => x"01",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"ff",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"fc",
           163 => x"10",
           164 => x"06",
           165 => x"92",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"fb",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"e7",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b5",
           272 => x"0b",
           273 => x"0b",
           274 => x"d5",
           275 => x"0b",
           276 => x"0b",
           277 => x"f5",
           278 => x"0b",
           279 => x"0b",
           280 => x"95",
           281 => x"0b",
           282 => x"0b",
           283 => x"b5",
           284 => x"0b",
           285 => x"0b",
           286 => x"d5",
           287 => x"0b",
           288 => x"0b",
           289 => x"f5",
           290 => x"0b",
           291 => x"0b",
           292 => x"93",
           293 => x"0b",
           294 => x"0b",
           295 => x"b2",
           296 => x"0b",
           297 => x"0b",
           298 => x"d2",
           299 => x"0b",
           300 => x"0b",
           301 => x"f2",
           302 => x"0b",
           303 => x"0b",
           304 => x"92",
           305 => x"0b",
           306 => x"0b",
           307 => x"b2",
           308 => x"0b",
           309 => x"0b",
           310 => x"d2",
           311 => x"0b",
           312 => x"0b",
           313 => x"f2",
           314 => x"0b",
           315 => x"0b",
           316 => x"92",
           317 => x"0b",
           318 => x"0b",
           319 => x"b2",
           320 => x"0b",
           321 => x"0b",
           322 => x"d2",
           323 => x"0b",
           324 => x"0b",
           325 => x"f2",
           326 => x"0b",
           327 => x"0b",
           328 => x"92",
           329 => x"0b",
           330 => x"0b",
           331 => x"b2",
           332 => x"0b",
           333 => x"0b",
           334 => x"d2",
           335 => x"0b",
           336 => x"0b",
           337 => x"f2",
           338 => x"0b",
           339 => x"0b",
           340 => x"91",
           341 => x"0b",
           342 => x"0b",
           343 => x"b0",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"2d",
           392 => x"08",
           393 => x"04",
           394 => x"0c",
           395 => x"2d",
           396 => x"08",
           397 => x"04",
           398 => x"0c",
           399 => x"2d",
           400 => x"08",
           401 => x"04",
           402 => x"0c",
           403 => x"2d",
           404 => x"08",
           405 => x"04",
           406 => x"0c",
           407 => x"2d",
           408 => x"08",
           409 => x"04",
           410 => x"0c",
           411 => x"2d",
           412 => x"08",
           413 => x"04",
           414 => x"0c",
           415 => x"2d",
           416 => x"08",
           417 => x"04",
           418 => x"0c",
           419 => x"2d",
           420 => x"08",
           421 => x"04",
           422 => x"0c",
           423 => x"2d",
           424 => x"08",
           425 => x"04",
           426 => x"0c",
           427 => x"2d",
           428 => x"08",
           429 => x"04",
           430 => x"0c",
           431 => x"2d",
           432 => x"08",
           433 => x"04",
           434 => x"0c",
           435 => x"2d",
           436 => x"08",
           437 => x"04",
           438 => x"0c",
           439 => x"2d",
           440 => x"08",
           441 => x"04",
           442 => x"0c",
           443 => x"2d",
           444 => x"08",
           445 => x"04",
           446 => x"0c",
           447 => x"82",
           448 => x"82",
           449 => x"82",
           450 => x"bd",
           451 => x"85",
           452 => x"a0",
           453 => x"85",
           454 => x"f0",
           455 => x"f8",
           456 => x"90",
           457 => x"f8",
           458 => x"bc",
           459 => x"f8",
           460 => x"90",
           461 => x"f8",
           462 => x"af",
           463 => x"f8",
           464 => x"90",
           465 => x"f8",
           466 => x"a3",
           467 => x"f8",
           468 => x"90",
           469 => x"f8",
           470 => x"a0",
           471 => x"f8",
           472 => x"90",
           473 => x"f8",
           474 => x"bd",
           475 => x"f8",
           476 => x"90",
           477 => x"f8",
           478 => x"a8",
           479 => x"f8",
           480 => x"90",
           481 => x"f8",
           482 => x"91",
           483 => x"f8",
           484 => x"90",
           485 => x"f8",
           486 => x"de",
           487 => x"f8",
           488 => x"90",
           489 => x"f8",
           490 => x"fd",
           491 => x"f8",
           492 => x"90",
           493 => x"f8",
           494 => x"9c",
           495 => x"f8",
           496 => x"90",
           497 => x"f8",
           498 => x"91",
           499 => x"f8",
           500 => x"90",
           501 => x"f8",
           502 => x"f5",
           503 => x"f8",
           504 => x"90",
           505 => x"f8",
           506 => x"e5",
           507 => x"f8",
           508 => x"90",
           509 => x"f8",
           510 => x"a2",
           511 => x"f8",
           512 => x"90",
           513 => x"f8",
           514 => x"e5",
           515 => x"f8",
           516 => x"90",
           517 => x"f8",
           518 => x"e6",
           519 => x"f8",
           520 => x"90",
           521 => x"f8",
           522 => x"8f",
           523 => x"f8",
           524 => x"90",
           525 => x"f8",
           526 => x"e8",
           527 => x"f8",
           528 => x"90",
           529 => x"f8",
           530 => x"93",
           531 => x"f8",
           532 => x"90",
           533 => x"f8",
           534 => x"f9",
           535 => x"f8",
           536 => x"90",
           537 => x"f8",
           538 => x"d7",
           539 => x"f8",
           540 => x"90",
           541 => x"f8",
           542 => x"e5",
           543 => x"f8",
           544 => x"90",
           545 => x"f8",
           546 => x"a7",
           547 => x"f8",
           548 => x"90",
           549 => x"f8",
           550 => x"db",
           551 => x"f8",
           552 => x"90",
           553 => x"f8",
           554 => x"95",
           555 => x"f8",
           556 => x"90",
           557 => x"f8",
           558 => x"d9",
           559 => x"f8",
           560 => x"90",
           561 => x"f8",
           562 => x"c0",
           563 => x"f8",
           564 => x"90",
           565 => x"f8",
           566 => x"e8",
           567 => x"f8",
           568 => x"90",
           569 => x"f8",
           570 => x"d2",
           571 => x"f8",
           572 => x"90",
           573 => x"f8",
           574 => x"b6",
           575 => x"f8",
           576 => x"90",
           577 => x"f8",
           578 => x"2d",
           579 => x"08",
           580 => x"04",
           581 => x"0c",
           582 => x"82",
           583 => x"82",
           584 => x"82",
           585 => x"80",
           586 => x"82",
           587 => x"82",
           588 => x"82",
           589 => x"a1",
           590 => x"85",
           591 => x"a0",
           592 => x"04",
           593 => x"10",
           594 => x"10",
           595 => x"10",
           596 => x"10",
           597 => x"10",
           598 => x"10",
           599 => x"10",
           600 => x"10",
           601 => x"04",
           602 => x"81",
           603 => x"83",
           604 => x"05",
           605 => x"10",
           606 => x"72",
           607 => x"51",
           608 => x"72",
           609 => x"06",
           610 => x"72",
           611 => x"10",
           612 => x"10",
           613 => x"ed",
           614 => x"53",
           615 => x"85",
           616 => x"9d",
           617 => x"38",
           618 => x"84",
           619 => x"0b",
           620 => x"9e",
           621 => x"51",
           622 => x"00",
           623 => x"08",
           624 => x"f8",
           625 => x"0d",
           626 => x"08",
           627 => x"82",
           628 => x"fc",
           629 => x"85",
           630 => x"05",
           631 => x"33",
           632 => x"08",
           633 => x"81",
           634 => x"f8",
           635 => x"0c",
           636 => x"06",
           637 => x"80",
           638 => x"da",
           639 => x"f8",
           640 => x"08",
           641 => x"85",
           642 => x"05",
           643 => x"f8",
           644 => x"08",
           645 => x"08",
           646 => x"31",
           647 => x"ec",
           648 => x"3d",
           649 => x"f8",
           650 => x"85",
           651 => x"82",
           652 => x"fe",
           653 => x"85",
           654 => x"05",
           655 => x"f8",
           656 => x"0c",
           657 => x"08",
           658 => x"52",
           659 => x"85",
           660 => x"05",
           661 => x"82",
           662 => x"8c",
           663 => x"85",
           664 => x"05",
           665 => x"70",
           666 => x"85",
           667 => x"05",
           668 => x"82",
           669 => x"fc",
           670 => x"81",
           671 => x"70",
           672 => x"38",
           673 => x"82",
           674 => x"88",
           675 => x"82",
           676 => x"51",
           677 => x"82",
           678 => x"04",
           679 => x"08",
           680 => x"f8",
           681 => x"0d",
           682 => x"08",
           683 => x"82",
           684 => x"fc",
           685 => x"85",
           686 => x"05",
           687 => x"f8",
           688 => x"0c",
           689 => x"08",
           690 => x"80",
           691 => x"38",
           692 => x"08",
           693 => x"81",
           694 => x"f8",
           695 => x"0c",
           696 => x"08",
           697 => x"ff",
           698 => x"f8",
           699 => x"0c",
           700 => x"08",
           701 => x"80",
           702 => x"82",
           703 => x"f8",
           704 => x"70",
           705 => x"f8",
           706 => x"08",
           707 => x"85",
           708 => x"05",
           709 => x"f8",
           710 => x"08",
           711 => x"71",
           712 => x"f8",
           713 => x"08",
           714 => x"85",
           715 => x"05",
           716 => x"39",
           717 => x"08",
           718 => x"70",
           719 => x"0c",
           720 => x"0d",
           721 => x"0c",
           722 => x"f8",
           723 => x"85",
           724 => x"3d",
           725 => x"f8",
           726 => x"08",
           727 => x"f4",
           728 => x"f8",
           729 => x"08",
           730 => x"82",
           731 => x"8c",
           732 => x"05",
           733 => x"08",
           734 => x"82",
           735 => x"88",
           736 => x"33",
           737 => x"06",
           738 => x"51",
           739 => x"84",
           740 => x"39",
           741 => x"08",
           742 => x"52",
           743 => x"85",
           744 => x"05",
           745 => x"82",
           746 => x"88",
           747 => x"81",
           748 => x"51",
           749 => x"80",
           750 => x"f8",
           751 => x"0c",
           752 => x"82",
           753 => x"90",
           754 => x"05",
           755 => x"08",
           756 => x"82",
           757 => x"90",
           758 => x"2e",
           759 => x"81",
           760 => x"f8",
           761 => x"08",
           762 => x"e8",
           763 => x"f8",
           764 => x"08",
           765 => x"53",
           766 => x"ff",
           767 => x"f8",
           768 => x"0c",
           769 => x"82",
           770 => x"8c",
           771 => x"05",
           772 => x"08",
           773 => x"82",
           774 => x"8c",
           775 => x"33",
           776 => x"8c",
           777 => x"82",
           778 => x"fc",
           779 => x"39",
           780 => x"08",
           781 => x"70",
           782 => x"f8",
           783 => x"08",
           784 => x"71",
           785 => x"85",
           786 => x"05",
           787 => x"52",
           788 => x"39",
           789 => x"85",
           790 => x"05",
           791 => x"f8",
           792 => x"08",
           793 => x"0c",
           794 => x"82",
           795 => x"04",
           796 => x"08",
           797 => x"f8",
           798 => x"0d",
           799 => x"08",
           800 => x"82",
           801 => x"fc",
           802 => x"85",
           803 => x"05",
           804 => x"80",
           805 => x"85",
           806 => x"05",
           807 => x"82",
           808 => x"90",
           809 => x"85",
           810 => x"05",
           811 => x"82",
           812 => x"90",
           813 => x"85",
           814 => x"05",
           815 => x"a9",
           816 => x"f8",
           817 => x"08",
           818 => x"85",
           819 => x"05",
           820 => x"71",
           821 => x"85",
           822 => x"05",
           823 => x"82",
           824 => x"fc",
           825 => x"be",
           826 => x"f8",
           827 => x"08",
           828 => x"ec",
           829 => x"3d",
           830 => x"f8",
           831 => x"85",
           832 => x"82",
           833 => x"f9",
           834 => x"0b",
           835 => x"08",
           836 => x"82",
           837 => x"88",
           838 => x"25",
           839 => x"85",
           840 => x"05",
           841 => x"85",
           842 => x"05",
           843 => x"82",
           844 => x"f4",
           845 => x"85",
           846 => x"05",
           847 => x"81",
           848 => x"f8",
           849 => x"0c",
           850 => x"08",
           851 => x"82",
           852 => x"fc",
           853 => x"85",
           854 => x"05",
           855 => x"b9",
           856 => x"f8",
           857 => x"08",
           858 => x"f8",
           859 => x"0c",
           860 => x"85",
           861 => x"05",
           862 => x"f8",
           863 => x"08",
           864 => x"0b",
           865 => x"08",
           866 => x"82",
           867 => x"f0",
           868 => x"85",
           869 => x"05",
           870 => x"82",
           871 => x"8c",
           872 => x"82",
           873 => x"88",
           874 => x"83",
           875 => x"85",
           876 => x"82",
           877 => x"f8",
           878 => x"82",
           879 => x"fc",
           880 => x"2e",
           881 => x"85",
           882 => x"05",
           883 => x"85",
           884 => x"05",
           885 => x"f8",
           886 => x"08",
           887 => x"ec",
           888 => x"3d",
           889 => x"f8",
           890 => x"85",
           891 => x"82",
           892 => x"fb",
           893 => x"0b",
           894 => x"08",
           895 => x"82",
           896 => x"88",
           897 => x"25",
           898 => x"85",
           899 => x"05",
           900 => x"85",
           901 => x"05",
           902 => x"82",
           903 => x"fc",
           904 => x"85",
           905 => x"05",
           906 => x"90",
           907 => x"f8",
           908 => x"08",
           909 => x"f8",
           910 => x"0c",
           911 => x"85",
           912 => x"05",
           913 => x"85",
           914 => x"05",
           915 => x"a2",
           916 => x"ec",
           917 => x"85",
           918 => x"05",
           919 => x"85",
           920 => x"05",
           921 => x"90",
           922 => x"f8",
           923 => x"08",
           924 => x"f8",
           925 => x"0c",
           926 => x"08",
           927 => x"70",
           928 => x"0c",
           929 => x"0d",
           930 => x"0c",
           931 => x"f8",
           932 => x"85",
           933 => x"3d",
           934 => x"82",
           935 => x"fc",
           936 => x"85",
           937 => x"05",
           938 => x"ff",
           939 => x"70",
           940 => x"08",
           941 => x"06",
           942 => x"08",
           943 => x"11",
           944 => x"08",
           945 => x"82",
           946 => x"88",
           947 => x"2a",
           948 => x"08",
           949 => x"82",
           950 => x"8c",
           951 => x"82",
           952 => x"8c",
           953 => x"51",
           954 => x"85",
           955 => x"05",
           956 => x"84",
           957 => x"39",
           958 => x"08",
           959 => x"70",
           960 => x"0c",
           961 => x"0d",
           962 => x"0c",
           963 => x"f8",
           964 => x"85",
           965 => x"3d",
           966 => x"82",
           967 => x"8c",
           968 => x"82",
           969 => x"88",
           970 => x"80",
           971 => x"85",
           972 => x"82",
           973 => x"54",
           974 => x"82",
           975 => x"04",
           976 => x"08",
           977 => x"f8",
           978 => x"0d",
           979 => x"85",
           980 => x"05",
           981 => x"85",
           982 => x"05",
           983 => x"3f",
           984 => x"08",
           985 => x"ec",
           986 => x"3d",
           987 => x"f8",
           988 => x"85",
           989 => x"82",
           990 => x"fd",
           991 => x"0b",
           992 => x"08",
           993 => x"80",
           994 => x"f8",
           995 => x"0c",
           996 => x"08",
           997 => x"82",
           998 => x"88",
           999 => x"b9",
          1000 => x"f8",
          1001 => x"08",
          1002 => x"38",
          1003 => x"85",
          1004 => x"05",
          1005 => x"38",
          1006 => x"08",
          1007 => x"10",
          1008 => x"08",
          1009 => x"82",
          1010 => x"fc",
          1011 => x"82",
          1012 => x"fc",
          1013 => x"b8",
          1014 => x"f8",
          1015 => x"08",
          1016 => x"e1",
          1017 => x"f8",
          1018 => x"08",
          1019 => x"08",
          1020 => x"26",
          1021 => x"85",
          1022 => x"05",
          1023 => x"f8",
          1024 => x"08",
          1025 => x"f8",
          1026 => x"0c",
          1027 => x"08",
          1028 => x"82",
          1029 => x"fc",
          1030 => x"82",
          1031 => x"f8",
          1032 => x"85",
          1033 => x"05",
          1034 => x"82",
          1035 => x"fc",
          1036 => x"85",
          1037 => x"05",
          1038 => x"82",
          1039 => x"8c",
          1040 => x"95",
          1041 => x"f8",
          1042 => x"08",
          1043 => x"38",
          1044 => x"08",
          1045 => x"70",
          1046 => x"08",
          1047 => x"51",
          1048 => x"85",
          1049 => x"05",
          1050 => x"85",
          1051 => x"05",
          1052 => x"85",
          1053 => x"05",
          1054 => x"ec",
          1055 => x"0d",
          1056 => x"0c",
          1057 => x"0d",
          1058 => x"70",
          1059 => x"74",
          1060 => x"e3",
          1061 => x"75",
          1062 => x"a0",
          1063 => x"ec",
          1064 => x"0c",
          1065 => x"54",
          1066 => x"74",
          1067 => x"a0",
          1068 => x"06",
          1069 => x"15",
          1070 => x"80",
          1071 => x"2b",
          1072 => x"05",
          1073 => x"56",
          1074 => x"82",
          1075 => x"53",
          1076 => x"08",
          1077 => x"3f",
          1078 => x"08",
          1079 => x"16",
          1080 => x"81",
          1081 => x"38",
          1082 => x"81",
          1083 => x"54",
          1084 => x"c9",
          1085 => x"73",
          1086 => x"0c",
          1087 => x"04",
          1088 => x"73",
          1089 => x"26",
          1090 => x"71",
          1091 => x"81",
          1092 => x"08",
          1093 => x"f4",
          1094 => x"39",
          1095 => x"51",
          1096 => x"81",
          1097 => x"80",
          1098 => x"eb",
          1099 => x"eb",
          1100 => x"b8",
          1101 => x"39",
          1102 => x"51",
          1103 => x"81",
          1104 => x"80",
          1105 => x"eb",
          1106 => x"cf",
          1107 => x"84",
          1108 => x"39",
          1109 => x"51",
          1110 => x"81",
          1111 => x"bb",
          1112 => x"d0",
          1113 => x"81",
          1114 => x"af",
          1115 => x"90",
          1116 => x"81",
          1117 => x"a3",
          1118 => x"c4",
          1119 => x"81",
          1120 => x"97",
          1121 => x"f0",
          1122 => x"81",
          1123 => x"8b",
          1124 => x"a0",
          1125 => x"81",
          1126 => x"ab",
          1127 => x"3d",
          1128 => x"3d",
          1129 => x"56",
          1130 => x"e7",
          1131 => x"87",
          1132 => x"51",
          1133 => x"74",
          1134 => x"ec",
          1135 => x"39",
          1136 => x"74",
          1137 => x"3f",
          1138 => x"08",
          1139 => x"fa",
          1140 => x"85",
          1141 => x"79",
          1142 => x"81",
          1143 => x"b0",
          1144 => x"3d",
          1145 => x"3d",
          1146 => x"84",
          1147 => x"05",
          1148 => x"80",
          1149 => x"81",
          1150 => x"07",
          1151 => x"57",
          1152 => x"56",
          1153 => x"26",
          1154 => x"56",
          1155 => x"70",
          1156 => x"51",
          1157 => x"74",
          1158 => x"81",
          1159 => x"8c",
          1160 => x"56",
          1161 => x"3f",
          1162 => x"08",
          1163 => x"ec",
          1164 => x"82",
          1165 => x"87",
          1166 => x"0c",
          1167 => x"08",
          1168 => x"d4",
          1169 => x"80",
          1170 => x"75",
          1171 => x"d6",
          1172 => x"ec",
          1173 => x"85",
          1174 => x"38",
          1175 => x"80",
          1176 => x"74",
          1177 => x"59",
          1178 => x"96",
          1179 => x"51",
          1180 => x"3f",
          1181 => x"05",
          1182 => x"80",
          1183 => x"81",
          1184 => x"2a",
          1185 => x"57",
          1186 => x"80",
          1187 => x"81",
          1188 => x"87",
          1189 => x"08",
          1190 => x"fe",
          1191 => x"56",
          1192 => x"ec",
          1193 => x"0d",
          1194 => x"0d",
          1195 => x"05",
          1196 => x"57",
          1197 => x"80",
          1198 => x"79",
          1199 => x"3f",
          1200 => x"08",
          1201 => x"80",
          1202 => x"75",
          1203 => x"38",
          1204 => x"55",
          1205 => x"85",
          1206 => x"52",
          1207 => x"2d",
          1208 => x"08",
          1209 => x"77",
          1210 => x"85",
          1211 => x"3d",
          1212 => x"3d",
          1213 => x"63",
          1214 => x"80",
          1215 => x"73",
          1216 => x"41",
          1217 => x"5e",
          1218 => x"52",
          1219 => x"51",
          1220 => x"81",
          1221 => x"a8",
          1222 => x"55",
          1223 => x"80",
          1224 => x"90",
          1225 => x"7b",
          1226 => x"38",
          1227 => x"74",
          1228 => x"7a",
          1229 => x"72",
          1230 => x"ee",
          1231 => x"9e",
          1232 => x"81",
          1233 => x"a8",
          1234 => x"15",
          1235 => x"74",
          1236 => x"7a",
          1237 => x"72",
          1238 => x"ee",
          1239 => x"fe",
          1240 => x"81",
          1241 => x"a8",
          1242 => x"15",
          1243 => x"74",
          1244 => x"7a",
          1245 => x"72",
          1246 => x"ef",
          1247 => x"de",
          1248 => x"81",
          1249 => x"a7",
          1250 => x"15",
          1251 => x"a7",
          1252 => x"88",
          1253 => x"94",
          1254 => x"3f",
          1255 => x"79",
          1256 => x"74",
          1257 => x"55",
          1258 => x"72",
          1259 => x"38",
          1260 => x"53",
          1261 => x"83",
          1262 => x"75",
          1263 => x"81",
          1264 => x"53",
          1265 => x"8b",
          1266 => x"fe",
          1267 => x"73",
          1268 => x"a0",
          1269 => x"3f",
          1270 => x"c2",
          1271 => x"98",
          1272 => x"3f",
          1273 => x"1c",
          1274 => x"fb",
          1275 => x"ec",
          1276 => x"70",
          1277 => x"57",
          1278 => x"09",
          1279 => x"38",
          1280 => x"82",
          1281 => x"98",
          1282 => x"2c",
          1283 => x"70",
          1284 => x"72",
          1285 => x"09",
          1286 => x"72",
          1287 => x"07",
          1288 => x"58",
          1289 => x"57",
          1290 => x"d4",
          1291 => x"2e",
          1292 => x"85",
          1293 => x"8c",
          1294 => x"53",
          1295 => x"fd",
          1296 => x"53",
          1297 => x"ec",
          1298 => x"0d",
          1299 => x"0d",
          1300 => x"33",
          1301 => x"53",
          1302 => x"52",
          1303 => x"3f",
          1304 => x"22",
          1305 => x"3f",
          1306 => x"54",
          1307 => x"53",
          1308 => x"33",
          1309 => x"c0",
          1310 => x"3f",
          1311 => x"84",
          1312 => x"3f",
          1313 => x"04",
          1314 => x"87",
          1315 => x"08",
          1316 => x"3f",
          1317 => x"eb",
          1318 => x"dc",
          1319 => x"3f",
          1320 => x"df",
          1321 => x"2a",
          1322 => x"51",
          1323 => x"2e",
          1324 => x"51",
          1325 => x"81",
          1326 => x"98",
          1327 => x"51",
          1328 => x"72",
          1329 => x"81",
          1330 => x"71",
          1331 => x"38",
          1332 => x"af",
          1333 => x"88",
          1334 => x"3f",
          1335 => x"a3",
          1336 => x"2a",
          1337 => x"51",
          1338 => x"2e",
          1339 => x"51",
          1340 => x"81",
          1341 => x"98",
          1342 => x"51",
          1343 => x"72",
          1344 => x"81",
          1345 => x"71",
          1346 => x"38",
          1347 => x"f3",
          1348 => x"ac",
          1349 => x"3f",
          1350 => x"e7",
          1351 => x"2a",
          1352 => x"51",
          1353 => x"2e",
          1354 => x"51",
          1355 => x"81",
          1356 => x"97",
          1357 => x"51",
          1358 => x"72",
          1359 => x"81",
          1360 => x"71",
          1361 => x"38",
          1362 => x"b7",
          1363 => x"d4",
          1364 => x"3f",
          1365 => x"ab",
          1366 => x"2a",
          1367 => x"51",
          1368 => x"2e",
          1369 => x"51",
          1370 => x"81",
          1371 => x"97",
          1372 => x"51",
          1373 => x"72",
          1374 => x"81",
          1375 => x"71",
          1376 => x"38",
          1377 => x"fb",
          1378 => x"fc",
          1379 => x"3f",
          1380 => x"ef",
          1381 => x"3f",
          1382 => x"04",
          1383 => x"77",
          1384 => x"a3",
          1385 => x"55",
          1386 => x"52",
          1387 => x"c0",
          1388 => x"82",
          1389 => x"54",
          1390 => x"81",
          1391 => x"bc",
          1392 => x"cc",
          1393 => x"f7",
          1394 => x"ec",
          1395 => x"05",
          1396 => x"ec",
          1397 => x"25",
          1398 => x"51",
          1399 => x"0b",
          1400 => x"e8",
          1401 => x"82",
          1402 => x"54",
          1403 => x"09",
          1404 => x"38",
          1405 => x"53",
          1406 => x"51",
          1407 => x"3f",
          1408 => x"08",
          1409 => x"38",
          1410 => x"08",
          1411 => x"3f",
          1412 => x"9c",
          1413 => x"8b",
          1414 => x"0b",
          1415 => x"80",
          1416 => x"0b",
          1417 => x"33",
          1418 => x"2e",
          1419 => x"8c",
          1420 => x"cc",
          1421 => x"75",
          1422 => x"3f",
          1423 => x"85",
          1424 => x"3d",
          1425 => x"3d",
          1426 => x"71",
          1427 => x"0c",
          1428 => x"52",
          1429 => x"cd",
          1430 => x"85",
          1431 => x"ff",
          1432 => x"7d",
          1433 => x"06",
          1434 => x"f1",
          1435 => x"3d",
          1436 => x"a7",
          1437 => x"53",
          1438 => x"86",
          1439 => x"fc",
          1440 => x"85",
          1441 => x"2e",
          1442 => x"f1",
          1443 => x"8a",
          1444 => x"5f",
          1445 => x"90",
          1446 => x"3f",
          1447 => x"46",
          1448 => x"52",
          1449 => x"f4",
          1450 => x"ff",
          1451 => x"f3",
          1452 => x"85",
          1453 => x"2b",
          1454 => x"51",
          1455 => x"c2",
          1456 => x"38",
          1457 => x"24",
          1458 => x"bd",
          1459 => x"38",
          1460 => x"90",
          1461 => x"2e",
          1462 => x"78",
          1463 => x"da",
          1464 => x"39",
          1465 => x"2e",
          1466 => x"78",
          1467 => x"85",
          1468 => x"bf",
          1469 => x"38",
          1470 => x"78",
          1471 => x"89",
          1472 => x"80",
          1473 => x"38",
          1474 => x"2e",
          1475 => x"78",
          1476 => x"89",
          1477 => x"86",
          1478 => x"83",
          1479 => x"38",
          1480 => x"24",
          1481 => x"81",
          1482 => x"d3",
          1483 => x"39",
          1484 => x"2e",
          1485 => x"89",
          1486 => x"3d",
          1487 => x"53",
          1488 => x"51",
          1489 => x"82",
          1490 => x"80",
          1491 => x"38",
          1492 => x"fc",
          1493 => x"84",
          1494 => x"fa",
          1495 => x"ec",
          1496 => x"fe",
          1497 => x"3d",
          1498 => x"53",
          1499 => x"51",
          1500 => x"82",
          1501 => x"86",
          1502 => x"ec",
          1503 => x"f2",
          1504 => x"ea",
          1505 => x"5c",
          1506 => x"27",
          1507 => x"61",
          1508 => x"70",
          1509 => x"0c",
          1510 => x"f5",
          1511 => x"39",
          1512 => x"80",
          1513 => x"84",
          1514 => x"aa",
          1515 => x"ec",
          1516 => x"fd",
          1517 => x"3d",
          1518 => x"53",
          1519 => x"51",
          1520 => x"82",
          1521 => x"80",
          1522 => x"38",
          1523 => x"f8",
          1524 => x"84",
          1525 => x"fe",
          1526 => x"ec",
          1527 => x"fd",
          1528 => x"f2",
          1529 => x"86",
          1530 => x"79",
          1531 => x"87",
          1532 => x"79",
          1533 => x"5b",
          1534 => x"61",
          1535 => x"eb",
          1536 => x"ff",
          1537 => x"ff",
          1538 => x"a6",
          1539 => x"85",
          1540 => x"2e",
          1541 => x"b4",
          1542 => x"11",
          1543 => x"05",
          1544 => x"3f",
          1545 => x"08",
          1546 => x"e9",
          1547 => x"fe",
          1548 => x"ff",
          1549 => x"a6",
          1550 => x"85",
          1551 => x"2e",
          1552 => x"81",
          1553 => x"9e",
          1554 => x"5a",
          1555 => x"a7",
          1556 => x"33",
          1557 => x"5a",
          1558 => x"2e",
          1559 => x"55",
          1560 => x"33",
          1561 => x"81",
          1562 => x"a3",
          1563 => x"1a",
          1564 => x"43",
          1565 => x"81",
          1566 => x"82",
          1567 => x"3d",
          1568 => x"53",
          1569 => x"51",
          1570 => x"82",
          1571 => x"80",
          1572 => x"84",
          1573 => x"78",
          1574 => x"38",
          1575 => x"08",
          1576 => x"39",
          1577 => x"33",
          1578 => x"2e",
          1579 => x"84",
          1580 => x"bc",
          1581 => x"da",
          1582 => x"80",
          1583 => x"82",
          1584 => x"44",
          1585 => x"84",
          1586 => x"78",
          1587 => x"38",
          1588 => x"08",
          1589 => x"82",
          1590 => x"59",
          1591 => x"88",
          1592 => x"b0",
          1593 => x"39",
          1594 => x"08",
          1595 => x"44",
          1596 => x"fc",
          1597 => x"84",
          1598 => x"da",
          1599 => x"ec",
          1600 => x"38",
          1601 => x"33",
          1602 => x"2e",
          1603 => x"84",
          1604 => x"80",
          1605 => x"84",
          1606 => x"78",
          1607 => x"38",
          1608 => x"08",
          1609 => x"82",
          1610 => x"59",
          1611 => x"88",
          1612 => x"a4",
          1613 => x"39",
          1614 => x"33",
          1615 => x"2e",
          1616 => x"84",
          1617 => x"99",
          1618 => x"d6",
          1619 => x"80",
          1620 => x"82",
          1621 => x"43",
          1622 => x"84",
          1623 => x"05",
          1624 => x"fe",
          1625 => x"ff",
          1626 => x"a3",
          1627 => x"85",
          1628 => x"2e",
          1629 => x"62",
          1630 => x"88",
          1631 => x"81",
          1632 => x"32",
          1633 => x"05",
          1634 => x"9f",
          1635 => x"06",
          1636 => x"5a",
          1637 => x"88",
          1638 => x"2e",
          1639 => x"42",
          1640 => x"51",
          1641 => x"a0",
          1642 => x"61",
          1643 => x"63",
          1644 => x"3f",
          1645 => x"51",
          1646 => x"f9",
          1647 => x"3d",
          1648 => x"53",
          1649 => x"51",
          1650 => x"82",
          1651 => x"80",
          1652 => x"38",
          1653 => x"fc",
          1654 => x"84",
          1655 => x"f6",
          1656 => x"ec",
          1657 => x"a4",
          1658 => x"02",
          1659 => x"33",
          1660 => x"81",
          1661 => x"3d",
          1662 => x"53",
          1663 => x"51",
          1664 => x"82",
          1665 => x"e1",
          1666 => x"39",
          1667 => x"54",
          1668 => x"f8",
          1669 => x"3f",
          1670 => x"79",
          1671 => x"3f",
          1672 => x"33",
          1673 => x"2e",
          1674 => x"9f",
          1675 => x"38",
          1676 => x"fc",
          1677 => x"84",
          1678 => x"9a",
          1679 => x"ec",
          1680 => x"91",
          1681 => x"02",
          1682 => x"33",
          1683 => x"81",
          1684 => x"b8",
          1685 => x"84",
          1686 => x"3f",
          1687 => x"b4",
          1688 => x"11",
          1689 => x"05",
          1690 => x"3f",
          1691 => x"08",
          1692 => x"a1",
          1693 => x"fe",
          1694 => x"ff",
          1695 => x"a3",
          1696 => x"85",
          1697 => x"2e",
          1698 => x"59",
          1699 => x"22",
          1700 => x"05",
          1701 => x"41",
          1702 => x"f0",
          1703 => x"84",
          1704 => x"ae",
          1705 => x"ec",
          1706 => x"f7",
          1707 => x"70",
          1708 => x"81",
          1709 => x"9f",
          1710 => x"f8",
          1711 => x"9f",
          1712 => x"45",
          1713 => x"78",
          1714 => x"c9",
          1715 => x"26",
          1716 => x"82",
          1717 => x"39",
          1718 => x"f0",
          1719 => x"84",
          1720 => x"ee",
          1721 => x"ec",
          1722 => x"92",
          1723 => x"02",
          1724 => x"79",
          1725 => x"5b",
          1726 => x"ff",
          1727 => x"f3",
          1728 => x"ea",
          1729 => x"39",
          1730 => x"f4",
          1731 => x"84",
          1732 => x"be",
          1733 => x"ec",
          1734 => x"f6",
          1735 => x"3d",
          1736 => x"53",
          1737 => x"51",
          1738 => x"82",
          1739 => x"80",
          1740 => x"60",
          1741 => x"59",
          1742 => x"41",
          1743 => x"f0",
          1744 => x"84",
          1745 => x"8a",
          1746 => x"ec",
          1747 => x"f6",
          1748 => x"70",
          1749 => x"81",
          1750 => x"9e",
          1751 => x"f8",
          1752 => x"9e",
          1753 => x"45",
          1754 => x"78",
          1755 => x"a5",
          1756 => x"27",
          1757 => x"3d",
          1758 => x"53",
          1759 => x"51",
          1760 => x"82",
          1761 => x"80",
          1762 => x"60",
          1763 => x"59",
          1764 => x"41",
          1765 => x"81",
          1766 => x"97",
          1767 => x"b2",
          1768 => x"ff",
          1769 => x"ff",
          1770 => x"9f",
          1771 => x"85",
          1772 => x"2e",
          1773 => x"63",
          1774 => x"a4",
          1775 => x"3f",
          1776 => x"04",
          1777 => x"80",
          1778 => x"84",
          1779 => x"86",
          1780 => x"ec",
          1781 => x"f5",
          1782 => x"52",
          1783 => x"51",
          1784 => x"63",
          1785 => x"82",
          1786 => x"80",
          1787 => x"38",
          1788 => x"08",
          1789 => x"dc",
          1790 => x"3f",
          1791 => x"81",
          1792 => x"96",
          1793 => x"96",
          1794 => x"39",
          1795 => x"51",
          1796 => x"80",
          1797 => x"39",
          1798 => x"f4",
          1799 => x"45",
          1800 => x"78",
          1801 => x"ed",
          1802 => x"06",
          1803 => x"2e",
          1804 => x"b4",
          1805 => x"05",
          1806 => x"3f",
          1807 => x"08",
          1808 => x"7a",
          1809 => x"38",
          1810 => x"89",
          1811 => x"2e",
          1812 => x"ca",
          1813 => x"2e",
          1814 => x"c2",
          1815 => x"a8",
          1816 => x"81",
          1817 => x"80",
          1818 => x"b0",
          1819 => x"ff",
          1820 => x"9b",
          1821 => x"39",
          1822 => x"52",
          1823 => x"b0",
          1824 => x"f0",
          1825 => x"7b",
          1826 => x"ac",
          1827 => x"81",
          1828 => x"b4",
          1829 => x"05",
          1830 => x"3f",
          1831 => x"54",
          1832 => x"f4",
          1833 => x"3d",
          1834 => x"51",
          1835 => x"82",
          1836 => x"82",
          1837 => x"80",
          1838 => x"80",
          1839 => x"80",
          1840 => x"80",
          1841 => x"ff",
          1842 => x"eb",
          1843 => x"85",
          1844 => x"85",
          1845 => x"70",
          1846 => x"70",
          1847 => x"25",
          1848 => x"5f",
          1849 => x"83",
          1850 => x"81",
          1851 => x"06",
          1852 => x"2e",
          1853 => x"1b",
          1854 => x"06",
          1855 => x"fe",
          1856 => x"81",
          1857 => x"32",
          1858 => x"8a",
          1859 => x"2e",
          1860 => x"f3",
          1861 => x"f4",
          1862 => x"c2",
          1863 => x"39",
          1864 => x"80",
          1865 => x"fc",
          1866 => x"94",
          1867 => x"54",
          1868 => x"80",
          1869 => x"e3",
          1870 => x"85",
          1871 => x"2b",
          1872 => x"53",
          1873 => x"52",
          1874 => x"c1",
          1875 => x"85",
          1876 => x"75",
          1877 => x"94",
          1878 => x"54",
          1879 => x"80",
          1880 => x"e3",
          1881 => x"85",
          1882 => x"2b",
          1883 => x"53",
          1884 => x"52",
          1885 => x"95",
          1886 => x"85",
          1887 => x"75",
          1888 => x"83",
          1889 => x"94",
          1890 => x"80",
          1891 => x"c0",
          1892 => x"80",
          1893 => x"82",
          1894 => x"80",
          1895 => x"82",
          1896 => x"89",
          1897 => x"d7",
          1898 => x"e4",
          1899 => x"3f",
          1900 => x"51",
          1901 => x"a9",
          1902 => x"be",
          1903 => x"ed",
          1904 => x"82",
          1905 => x"fe",
          1906 => x"52",
          1907 => x"88",
          1908 => x"c4",
          1909 => x"ec",
          1910 => x"06",
          1911 => x"14",
          1912 => x"80",
          1913 => x"71",
          1914 => x"0c",
          1915 => x"04",
          1916 => x"76",
          1917 => x"55",
          1918 => x"54",
          1919 => x"81",
          1920 => x"33",
          1921 => x"2e",
          1922 => x"86",
          1923 => x"53",
          1924 => x"33",
          1925 => x"2e",
          1926 => x"86",
          1927 => x"53",
          1928 => x"52",
          1929 => x"09",
          1930 => x"38",
          1931 => x"12",
          1932 => x"33",
          1933 => x"a2",
          1934 => x"81",
          1935 => x"2e",
          1936 => x"ea",
          1937 => x"81",
          1938 => x"72",
          1939 => x"70",
          1940 => x"38",
          1941 => x"80",
          1942 => x"73",
          1943 => x"72",
          1944 => x"70",
          1945 => x"81",
          1946 => x"81",
          1947 => x"32",
          1948 => x"05",
          1949 => x"76",
          1950 => x"51",
          1951 => x"88",
          1952 => x"70",
          1953 => x"34",
          1954 => x"72",
          1955 => x"85",
          1956 => x"3d",
          1957 => x"3d",
          1958 => x"72",
          1959 => x"91",
          1960 => x"fc",
          1961 => x"51",
          1962 => x"82",
          1963 => x"85",
          1964 => x"83",
          1965 => x"72",
          1966 => x"0c",
          1967 => x"04",
          1968 => x"76",
          1969 => x"ff",
          1970 => x"81",
          1971 => x"26",
          1972 => x"83",
          1973 => x"05",
          1974 => x"70",
          1975 => x"8a",
          1976 => x"33",
          1977 => x"70",
          1978 => x"fe",
          1979 => x"33",
          1980 => x"70",
          1981 => x"f2",
          1982 => x"33",
          1983 => x"70",
          1984 => x"e6",
          1985 => x"22",
          1986 => x"74",
          1987 => x"80",
          1988 => x"13",
          1989 => x"52",
          1990 => x"26",
          1991 => x"81",
          1992 => x"98",
          1993 => x"22",
          1994 => x"bc",
          1995 => x"33",
          1996 => x"b8",
          1997 => x"33",
          1998 => x"b4",
          1999 => x"33",
          2000 => x"b0",
          2001 => x"33",
          2002 => x"ac",
          2003 => x"33",
          2004 => x"a8",
          2005 => x"c0",
          2006 => x"73",
          2007 => x"a0",
          2008 => x"87",
          2009 => x"0c",
          2010 => x"82",
          2011 => x"86",
          2012 => x"f3",
          2013 => x"5b",
          2014 => x"9c",
          2015 => x"0c",
          2016 => x"bc",
          2017 => x"7b",
          2018 => x"98",
          2019 => x"79",
          2020 => x"87",
          2021 => x"08",
          2022 => x"1c",
          2023 => x"98",
          2024 => x"79",
          2025 => x"87",
          2026 => x"08",
          2027 => x"1c",
          2028 => x"98",
          2029 => x"79",
          2030 => x"87",
          2031 => x"08",
          2032 => x"1c",
          2033 => x"98",
          2034 => x"79",
          2035 => x"80",
          2036 => x"83",
          2037 => x"59",
          2038 => x"ff",
          2039 => x"1b",
          2040 => x"1b",
          2041 => x"1b",
          2042 => x"1b",
          2043 => x"1b",
          2044 => x"83",
          2045 => x"52",
          2046 => x"51",
          2047 => x"8f",
          2048 => x"ff",
          2049 => x"8f",
          2050 => x"09",
          2051 => x"9f",
          2052 => x"52",
          2053 => x"8c",
          2054 => x"0d",
          2055 => x"0d",
          2056 => x"8c",
          2057 => x"ff",
          2058 => x"56",
          2059 => x"84",
          2060 => x"2e",
          2061 => x"c0",
          2062 => x"70",
          2063 => x"2a",
          2064 => x"53",
          2065 => x"80",
          2066 => x"71",
          2067 => x"81",
          2068 => x"70",
          2069 => x"81",
          2070 => x"06",
          2071 => x"80",
          2072 => x"71",
          2073 => x"81",
          2074 => x"70",
          2075 => x"73",
          2076 => x"51",
          2077 => x"80",
          2078 => x"2e",
          2079 => x"c0",
          2080 => x"75",
          2081 => x"82",
          2082 => x"87",
          2083 => x"fb",
          2084 => x"9f",
          2085 => x"84",
          2086 => x"81",
          2087 => x"55",
          2088 => x"94",
          2089 => x"80",
          2090 => x"87",
          2091 => x"51",
          2092 => x"96",
          2093 => x"06",
          2094 => x"70",
          2095 => x"38",
          2096 => x"70",
          2097 => x"51",
          2098 => x"72",
          2099 => x"81",
          2100 => x"70",
          2101 => x"38",
          2102 => x"70",
          2103 => x"51",
          2104 => x"38",
          2105 => x"06",
          2106 => x"94",
          2107 => x"80",
          2108 => x"87",
          2109 => x"52",
          2110 => x"87",
          2111 => x"f9",
          2112 => x"54",
          2113 => x"70",
          2114 => x"53",
          2115 => x"77",
          2116 => x"38",
          2117 => x"06",
          2118 => x"84",
          2119 => x"81",
          2120 => x"57",
          2121 => x"c0",
          2122 => x"75",
          2123 => x"38",
          2124 => x"94",
          2125 => x"70",
          2126 => x"81",
          2127 => x"52",
          2128 => x"8c",
          2129 => x"2a",
          2130 => x"51",
          2131 => x"38",
          2132 => x"70",
          2133 => x"51",
          2134 => x"8d",
          2135 => x"2a",
          2136 => x"51",
          2137 => x"be",
          2138 => x"ff",
          2139 => x"c0",
          2140 => x"70",
          2141 => x"38",
          2142 => x"90",
          2143 => x"0c",
          2144 => x"33",
          2145 => x"06",
          2146 => x"70",
          2147 => x"76",
          2148 => x"0c",
          2149 => x"04",
          2150 => x"82",
          2151 => x"70",
          2152 => x"54",
          2153 => x"94",
          2154 => x"80",
          2155 => x"87",
          2156 => x"51",
          2157 => x"82",
          2158 => x"06",
          2159 => x"70",
          2160 => x"38",
          2161 => x"06",
          2162 => x"94",
          2163 => x"80",
          2164 => x"87",
          2165 => x"52",
          2166 => x"81",
          2167 => x"85",
          2168 => x"84",
          2169 => x"fe",
          2170 => x"84",
          2171 => x"81",
          2172 => x"53",
          2173 => x"84",
          2174 => x"2e",
          2175 => x"c0",
          2176 => x"71",
          2177 => x"2a",
          2178 => x"51",
          2179 => x"52",
          2180 => x"a0",
          2181 => x"ff",
          2182 => x"c0",
          2183 => x"70",
          2184 => x"38",
          2185 => x"90",
          2186 => x"70",
          2187 => x"98",
          2188 => x"51",
          2189 => x"ec",
          2190 => x"0d",
          2191 => x"0d",
          2192 => x"80",
          2193 => x"2a",
          2194 => x"51",
          2195 => x"84",
          2196 => x"c0",
          2197 => x"82",
          2198 => x"87",
          2199 => x"08",
          2200 => x"0c",
          2201 => x"94",
          2202 => x"98",
          2203 => x"9e",
          2204 => x"84",
          2205 => x"c0",
          2206 => x"82",
          2207 => x"87",
          2208 => x"08",
          2209 => x"0c",
          2210 => x"ac",
          2211 => x"a8",
          2212 => x"9e",
          2213 => x"84",
          2214 => x"c0",
          2215 => x"82",
          2216 => x"87",
          2217 => x"08",
          2218 => x"0c",
          2219 => x"bc",
          2220 => x"b8",
          2221 => x"9e",
          2222 => x"84",
          2223 => x"c0",
          2224 => x"82",
          2225 => x"87",
          2226 => x"08",
          2227 => x"84",
          2228 => x"c0",
          2229 => x"82",
          2230 => x"87",
          2231 => x"08",
          2232 => x"0c",
          2233 => x"8c",
          2234 => x"d0",
          2235 => x"82",
          2236 => x"80",
          2237 => x"9e",
          2238 => x"84",
          2239 => x"51",
          2240 => x"80",
          2241 => x"81",
          2242 => x"84",
          2243 => x"0b",
          2244 => x"90",
          2245 => x"80",
          2246 => x"52",
          2247 => x"2e",
          2248 => x"52",
          2249 => x"d6",
          2250 => x"87",
          2251 => x"08",
          2252 => x"0a",
          2253 => x"52",
          2254 => x"83",
          2255 => x"71",
          2256 => x"34",
          2257 => x"c0",
          2258 => x"70",
          2259 => x"06",
          2260 => x"70",
          2261 => x"38",
          2262 => x"82",
          2263 => x"80",
          2264 => x"9e",
          2265 => x"a0",
          2266 => x"51",
          2267 => x"80",
          2268 => x"81",
          2269 => x"84",
          2270 => x"0b",
          2271 => x"90",
          2272 => x"80",
          2273 => x"52",
          2274 => x"2e",
          2275 => x"52",
          2276 => x"da",
          2277 => x"87",
          2278 => x"08",
          2279 => x"80",
          2280 => x"52",
          2281 => x"83",
          2282 => x"71",
          2283 => x"34",
          2284 => x"c0",
          2285 => x"70",
          2286 => x"06",
          2287 => x"70",
          2288 => x"38",
          2289 => x"82",
          2290 => x"80",
          2291 => x"9e",
          2292 => x"81",
          2293 => x"51",
          2294 => x"80",
          2295 => x"81",
          2296 => x"84",
          2297 => x"0b",
          2298 => x"90",
          2299 => x"c0",
          2300 => x"52",
          2301 => x"2e",
          2302 => x"52",
          2303 => x"de",
          2304 => x"87",
          2305 => x"08",
          2306 => x"06",
          2307 => x"70",
          2308 => x"38",
          2309 => x"82",
          2310 => x"87",
          2311 => x"08",
          2312 => x"06",
          2313 => x"51",
          2314 => x"82",
          2315 => x"80",
          2316 => x"9e",
          2317 => x"84",
          2318 => x"52",
          2319 => x"2e",
          2320 => x"52",
          2321 => x"e1",
          2322 => x"9e",
          2323 => x"83",
          2324 => x"84",
          2325 => x"51",
          2326 => x"e2",
          2327 => x"87",
          2328 => x"08",
          2329 => x"51",
          2330 => x"80",
          2331 => x"81",
          2332 => x"84",
          2333 => x"c0",
          2334 => x"70",
          2335 => x"51",
          2336 => x"e4",
          2337 => x"0d",
          2338 => x"0d",
          2339 => x"51",
          2340 => x"82",
          2341 => x"54",
          2342 => x"88",
          2343 => x"b4",
          2344 => x"3f",
          2345 => x"51",
          2346 => x"82",
          2347 => x"54",
          2348 => x"93",
          2349 => x"b0",
          2350 => x"b4",
          2351 => x"52",
          2352 => x"51",
          2353 => x"82",
          2354 => x"54",
          2355 => x"93",
          2356 => x"a8",
          2357 => x"ac",
          2358 => x"52",
          2359 => x"51",
          2360 => x"82",
          2361 => x"54",
          2362 => x"93",
          2363 => x"90",
          2364 => x"94",
          2365 => x"52",
          2366 => x"51",
          2367 => x"82",
          2368 => x"54",
          2369 => x"93",
          2370 => x"98",
          2371 => x"9c",
          2372 => x"52",
          2373 => x"51",
          2374 => x"82",
          2375 => x"54",
          2376 => x"93",
          2377 => x"a0",
          2378 => x"a4",
          2379 => x"52",
          2380 => x"51",
          2381 => x"82",
          2382 => x"54",
          2383 => x"8d",
          2384 => x"e0",
          2385 => x"f6",
          2386 => x"92",
          2387 => x"e3",
          2388 => x"80",
          2389 => x"82",
          2390 => x"52",
          2391 => x"51",
          2392 => x"82",
          2393 => x"54",
          2394 => x"8d",
          2395 => x"e2",
          2396 => x"f7",
          2397 => x"e6",
          2398 => x"d5",
          2399 => x"80",
          2400 => x"81",
          2401 => x"83",
          2402 => x"84",
          2403 => x"73",
          2404 => x"38",
          2405 => x"51",
          2406 => x"82",
          2407 => x"54",
          2408 => x"88",
          2409 => x"ec",
          2410 => x"3f",
          2411 => x"33",
          2412 => x"2e",
          2413 => x"f7",
          2414 => x"b2",
          2415 => x"de",
          2416 => x"80",
          2417 => x"81",
          2418 => x"83",
          2419 => x"f8",
          2420 => x"9a",
          2421 => x"b8",
          2422 => x"f8",
          2423 => x"fe",
          2424 => x"bc",
          2425 => x"f8",
          2426 => x"f2",
          2427 => x"c0",
          2428 => x"f8",
          2429 => x"e6",
          2430 => x"94",
          2431 => x"3f",
          2432 => x"22",
          2433 => x"9c",
          2434 => x"3f",
          2435 => x"08",
          2436 => x"c0",
          2437 => x"d1",
          2438 => x"85",
          2439 => x"bd",
          2440 => x"82",
          2441 => x"51",
          2442 => x"74",
          2443 => x"08",
          2444 => x"52",
          2445 => x"51",
          2446 => x"82",
          2447 => x"54",
          2448 => x"b0",
          2449 => x"cc",
          2450 => x"84",
          2451 => x"51",
          2452 => x"82",
          2453 => x"54",
          2454 => x"52",
          2455 => x"08",
          2456 => x"3f",
          2457 => x"ec",
          2458 => x"73",
          2459 => x"f0",
          2460 => x"3f",
          2461 => x"33",
          2462 => x"2e",
          2463 => x"84",
          2464 => x"bd",
          2465 => x"74",
          2466 => x"3f",
          2467 => x"08",
          2468 => x"c0",
          2469 => x"ec",
          2470 => x"f1",
          2471 => x"85",
          2472 => x"53",
          2473 => x"fa",
          2474 => x"b2",
          2475 => x"d8",
          2476 => x"3f",
          2477 => x"04",
          2478 => x"02",
          2479 => x"ff",
          2480 => x"84",
          2481 => x"71",
          2482 => x"81",
          2483 => x"08",
          2484 => x"c8",
          2485 => x"81",
          2486 => x"97",
          2487 => x"d8",
          2488 => x"81",
          2489 => x"8b",
          2490 => x"e4",
          2491 => x"81",
          2492 => x"80",
          2493 => x"3d",
          2494 => x"88",
          2495 => x"80",
          2496 => x"96",
          2497 => x"82",
          2498 => x"87",
          2499 => x"0c",
          2500 => x"0d",
          2501 => x"33",
          2502 => x"2e",
          2503 => x"85",
          2504 => x"ed",
          2505 => x"fc",
          2506 => x"80",
          2507 => x"72",
          2508 => x"9c",
          2509 => x"05",
          2510 => x"0c",
          2511 => x"9c",
          2512 => x"71",
          2513 => x"38",
          2514 => x"2d",
          2515 => x"04",
          2516 => x"02",
          2517 => x"82",
          2518 => x"76",
          2519 => x"0c",
          2520 => x"ad",
          2521 => x"9c",
          2522 => x"3d",
          2523 => x"3d",
          2524 => x"73",
          2525 => x"ff",
          2526 => x"71",
          2527 => x"38",
          2528 => x"06",
          2529 => x"54",
          2530 => x"e7",
          2531 => x"0d",
          2532 => x"0d",
          2533 => x"f4",
          2534 => x"9c",
          2535 => x"54",
          2536 => x"81",
          2537 => x"53",
          2538 => x"8e",
          2539 => x"ff",
          2540 => x"14",
          2541 => x"3f",
          2542 => x"82",
          2543 => x"86",
          2544 => x"ec",
          2545 => x"68",
          2546 => x"70",
          2547 => x"33",
          2548 => x"2e",
          2549 => x"75",
          2550 => x"81",
          2551 => x"38",
          2552 => x"70",
          2553 => x"33",
          2554 => x"75",
          2555 => x"81",
          2556 => x"81",
          2557 => x"75",
          2558 => x"81",
          2559 => x"82",
          2560 => x"81",
          2561 => x"56",
          2562 => x"09",
          2563 => x"38",
          2564 => x"71",
          2565 => x"81",
          2566 => x"59",
          2567 => x"9f",
          2568 => x"53",
          2569 => x"97",
          2570 => x"2b",
          2571 => x"11",
          2572 => x"7b",
          2573 => x"5d",
          2574 => x"51",
          2575 => x"75",
          2576 => x"70",
          2577 => x"70",
          2578 => x"25",
          2579 => x"32",
          2580 => x"05",
          2581 => x"80",
          2582 => x"53",
          2583 => x"55",
          2584 => x"2e",
          2585 => x"84",
          2586 => x"81",
          2587 => x"57",
          2588 => x"2e",
          2589 => x"75",
          2590 => x"76",
          2591 => x"e0",
          2592 => x"ff",
          2593 => x"73",
          2594 => x"81",
          2595 => x"80",
          2596 => x"38",
          2597 => x"2e",
          2598 => x"73",
          2599 => x"8b",
          2600 => x"c2",
          2601 => x"38",
          2602 => x"73",
          2603 => x"81",
          2604 => x"8f",
          2605 => x"d5",
          2606 => x"38",
          2607 => x"24",
          2608 => x"80",
          2609 => x"38",
          2610 => x"73",
          2611 => x"80",
          2612 => x"ef",
          2613 => x"19",
          2614 => x"59",
          2615 => x"33",
          2616 => x"75",
          2617 => x"81",
          2618 => x"70",
          2619 => x"55",
          2620 => x"79",
          2621 => x"90",
          2622 => x"16",
          2623 => x"7b",
          2624 => x"a0",
          2625 => x"3f",
          2626 => x"53",
          2627 => x"e9",
          2628 => x"fc",
          2629 => x"81",
          2630 => x"72",
          2631 => x"aa",
          2632 => x"fb",
          2633 => x"39",
          2634 => x"83",
          2635 => x"59",
          2636 => x"82",
          2637 => x"88",
          2638 => x"8a",
          2639 => x"90",
          2640 => x"75",
          2641 => x"3f",
          2642 => x"79",
          2643 => x"81",
          2644 => x"72",
          2645 => x"38",
          2646 => x"59",
          2647 => x"84",
          2648 => x"58",
          2649 => x"80",
          2650 => x"09",
          2651 => x"72",
          2652 => x"51",
          2653 => x"74",
          2654 => x"38",
          2655 => x"8a",
          2656 => x"81",
          2657 => x"07",
          2658 => x"0b",
          2659 => x"57",
          2660 => x"51",
          2661 => x"82",
          2662 => x"81",
          2663 => x"53",
          2664 => x"ca",
          2665 => x"85",
          2666 => x"89",
          2667 => x"38",
          2668 => x"75",
          2669 => x"84",
          2670 => x"53",
          2671 => x"06",
          2672 => x"53",
          2673 => x"81",
          2674 => x"81",
          2675 => x"81",
          2676 => x"07",
          2677 => x"54",
          2678 => x"26",
          2679 => x"ff",
          2680 => x"84",
          2681 => x"06",
          2682 => x"80",
          2683 => x"96",
          2684 => x"e0",
          2685 => x"73",
          2686 => x"57",
          2687 => x"06",
          2688 => x"54",
          2689 => x"a0",
          2690 => x"2a",
          2691 => x"54",
          2692 => x"38",
          2693 => x"76",
          2694 => x"38",
          2695 => x"f1",
          2696 => x"06",
          2697 => x"38",
          2698 => x"56",
          2699 => x"26",
          2700 => x"3d",
          2701 => x"05",
          2702 => x"ff",
          2703 => x"53",
          2704 => x"cd",
          2705 => x"38",
          2706 => x"56",
          2707 => x"27",
          2708 => x"a0",
          2709 => x"3f",
          2710 => x"3d",
          2711 => x"3d",
          2712 => x"70",
          2713 => x"52",
          2714 => x"73",
          2715 => x"3f",
          2716 => x"04",
          2717 => x"74",
          2718 => x"0c",
          2719 => x"05",
          2720 => x"fa",
          2721 => x"9c",
          2722 => x"80",
          2723 => x"0b",
          2724 => x"0c",
          2725 => x"04",
          2726 => x"82",
          2727 => x"76",
          2728 => x"0c",
          2729 => x"05",
          2730 => x"53",
          2731 => x"72",
          2732 => x"0c",
          2733 => x"04",
          2734 => x"77",
          2735 => x"f8",
          2736 => x"54",
          2737 => x"54",
          2738 => x"80",
          2739 => x"9c",
          2740 => x"71",
          2741 => x"ec",
          2742 => x"06",
          2743 => x"2e",
          2744 => x"72",
          2745 => x"38",
          2746 => x"70",
          2747 => x"70",
          2748 => x"51",
          2749 => x"2e",
          2750 => x"80",
          2751 => x"ff",
          2752 => x"39",
          2753 => x"c6",
          2754 => x"52",
          2755 => x"ff",
          2756 => x"14",
          2757 => x"34",
          2758 => x"72",
          2759 => x"3f",
          2760 => x"73",
          2761 => x"72",
          2762 => x"f7",
          2763 => x"53",
          2764 => x"ec",
          2765 => x"0d",
          2766 => x"0d",
          2767 => x"08",
          2768 => x"f8",
          2769 => x"76",
          2770 => x"ec",
          2771 => x"9c",
          2772 => x"3d",
          2773 => x"3d",
          2774 => x"5a",
          2775 => x"7a",
          2776 => x"08",
          2777 => x"53",
          2778 => x"09",
          2779 => x"38",
          2780 => x"0c",
          2781 => x"ad",
          2782 => x"06",
          2783 => x"76",
          2784 => x"0c",
          2785 => x"33",
          2786 => x"73",
          2787 => x"81",
          2788 => x"38",
          2789 => x"05",
          2790 => x"08",
          2791 => x"53",
          2792 => x"2e",
          2793 => x"57",
          2794 => x"2e",
          2795 => x"39",
          2796 => x"13",
          2797 => x"08",
          2798 => x"53",
          2799 => x"55",
          2800 => x"81",
          2801 => x"14",
          2802 => x"88",
          2803 => x"27",
          2804 => x"f5",
          2805 => x"53",
          2806 => x"89",
          2807 => x"38",
          2808 => x"55",
          2809 => x"8a",
          2810 => x"a0",
          2811 => x"ca",
          2812 => x"74",
          2813 => x"e0",
          2814 => x"ff",
          2815 => x"d0",
          2816 => x"ff",
          2817 => x"90",
          2818 => x"38",
          2819 => x"81",
          2820 => x"53",
          2821 => x"ca",
          2822 => x"27",
          2823 => x"52",
          2824 => x"e9",
          2825 => x"ec",
          2826 => x"08",
          2827 => x"0c",
          2828 => x"33",
          2829 => x"ff",
          2830 => x"80",
          2831 => x"74",
          2832 => x"55",
          2833 => x"81",
          2834 => x"85",
          2835 => x"3d",
          2836 => x"3d",
          2837 => x"5a",
          2838 => x"7a",
          2839 => x"08",
          2840 => x"53",
          2841 => x"09",
          2842 => x"38",
          2843 => x"0c",
          2844 => x"ad",
          2845 => x"06",
          2846 => x"76",
          2847 => x"0c",
          2848 => x"33",
          2849 => x"73",
          2850 => x"81",
          2851 => x"38",
          2852 => x"05",
          2853 => x"08",
          2854 => x"53",
          2855 => x"2e",
          2856 => x"57",
          2857 => x"2e",
          2858 => x"39",
          2859 => x"13",
          2860 => x"08",
          2861 => x"53",
          2862 => x"55",
          2863 => x"81",
          2864 => x"14",
          2865 => x"88",
          2866 => x"27",
          2867 => x"f5",
          2868 => x"53",
          2869 => x"89",
          2870 => x"38",
          2871 => x"55",
          2872 => x"8a",
          2873 => x"a0",
          2874 => x"ca",
          2875 => x"74",
          2876 => x"e0",
          2877 => x"ff",
          2878 => x"d0",
          2879 => x"ff",
          2880 => x"90",
          2881 => x"38",
          2882 => x"81",
          2883 => x"53",
          2884 => x"ca",
          2885 => x"27",
          2886 => x"52",
          2887 => x"ed",
          2888 => x"ec",
          2889 => x"08",
          2890 => x"0c",
          2891 => x"33",
          2892 => x"ff",
          2893 => x"80",
          2894 => x"74",
          2895 => x"55",
          2896 => x"81",
          2897 => x"85",
          2898 => x"3d",
          2899 => x"3d",
          2900 => x"2b",
          2901 => x"79",
          2902 => x"98",
          2903 => x"73",
          2904 => x"54",
          2905 => x"51",
          2906 => x"81",
          2907 => x"33",
          2908 => x"74",
          2909 => x"71",
          2910 => x"12",
          2911 => x"88",
          2912 => x"33",
          2913 => x"53",
          2914 => x"72",
          2915 => x"06",
          2916 => x"54",
          2917 => x"82",
          2918 => x"85",
          2919 => x"fc",
          2920 => x"02",
          2921 => x"05",
          2922 => x"54",
          2923 => x"80",
          2924 => x"88",
          2925 => x"3f",
          2926 => x"d5",
          2927 => x"f2",
          2928 => x"33",
          2929 => x"71",
          2930 => x"81",
          2931 => x"de",
          2932 => x"f3",
          2933 => x"73",
          2934 => x"0d",
          2935 => x"0d",
          2936 => x"05",
          2937 => x"02",
          2938 => x"05",
          2939 => x"c4",
          2940 => x"2b",
          2941 => x"11",
          2942 => x"59",
          2943 => x"74",
          2944 => x"38",
          2945 => x"87",
          2946 => x"c4",
          2947 => x"2b",
          2948 => x"11",
          2949 => x"55",
          2950 => x"5a",
          2951 => x"82",
          2952 => x"75",
          2953 => x"c4",
          2954 => x"2b",
          2955 => x"11",
          2956 => x"5a",
          2957 => x"a7",
          2958 => x"78",
          2959 => x"ff",
          2960 => x"82",
          2961 => x"81",
          2962 => x"82",
          2963 => x"74",
          2964 => x"55",
          2965 => x"87",
          2966 => x"82",
          2967 => x"77",
          2968 => x"38",
          2969 => x"08",
          2970 => x"2e",
          2971 => x"85",
          2972 => x"74",
          2973 => x"3d",
          2974 => x"76",
          2975 => x"75",
          2976 => x"9f",
          2977 => x"c0",
          2978 => x"51",
          2979 => x"3f",
          2980 => x"08",
          2981 => x"fc",
          2982 => x"0d",
          2983 => x"0d",
          2984 => x"53",
          2985 => x"08",
          2986 => x"2e",
          2987 => x"51",
          2988 => x"80",
          2989 => x"14",
          2990 => x"54",
          2991 => x"e6",
          2992 => x"82",
          2993 => x"82",
          2994 => x"52",
          2995 => x"95",
          2996 => x"80",
          2997 => x"82",
          2998 => x"51",
          2999 => x"80",
          3000 => x"c0",
          3001 => x"0d",
          3002 => x"0d",
          3003 => x"52",
          3004 => x"08",
          3005 => x"c8",
          3006 => x"ec",
          3007 => x"38",
          3008 => x"08",
          3009 => x"52",
          3010 => x"52",
          3011 => x"b3",
          3012 => x"ec",
          3013 => x"b9",
          3014 => x"ff",
          3015 => x"82",
          3016 => x"55",
          3017 => x"85",
          3018 => x"9c",
          3019 => x"ec",
          3020 => x"70",
          3021 => x"80",
          3022 => x"53",
          3023 => x"17",
          3024 => x"52",
          3025 => x"3f",
          3026 => x"09",
          3027 => x"b0",
          3028 => x"0d",
          3029 => x"0d",
          3030 => x"ad",
          3031 => x"5a",
          3032 => x"58",
          3033 => x"85",
          3034 => x"80",
          3035 => x"82",
          3036 => x"81",
          3037 => x"0b",
          3038 => x"08",
          3039 => x"f8",
          3040 => x"70",
          3041 => x"86",
          3042 => x"85",
          3043 => x"2e",
          3044 => x"51",
          3045 => x"3f",
          3046 => x"08",
          3047 => x"55",
          3048 => x"85",
          3049 => x"8e",
          3050 => x"ec",
          3051 => x"70",
          3052 => x"80",
          3053 => x"09",
          3054 => x"05",
          3055 => x"9f",
          3056 => x"55",
          3057 => x"85",
          3058 => x"aa",
          3059 => x"c0",
          3060 => x"08",
          3061 => x"dc",
          3062 => x"85",
          3063 => x"2e",
          3064 => x"fd",
          3065 => x"86",
          3066 => x"2e",
          3067 => x"9b",
          3068 => x"79",
          3069 => x"b2",
          3070 => x"ff",
          3071 => x"ab",
          3072 => x"82",
          3073 => x"74",
          3074 => x"77",
          3075 => x"0c",
          3076 => x"04",
          3077 => x"7c",
          3078 => x"71",
          3079 => x"59",
          3080 => x"a0",
          3081 => x"06",
          3082 => x"33",
          3083 => x"77",
          3084 => x"38",
          3085 => x"5b",
          3086 => x"56",
          3087 => x"a0",
          3088 => x"06",
          3089 => x"75",
          3090 => x"80",
          3091 => x"2b",
          3092 => x"11",
          3093 => x"51",
          3094 => x"e0",
          3095 => x"ec",
          3096 => x"52",
          3097 => x"ff",
          3098 => x"82",
          3099 => x"80",
          3100 => x"14",
          3101 => x"81",
          3102 => x"73",
          3103 => x"38",
          3104 => x"e5",
          3105 => x"81",
          3106 => x"3d",
          3107 => x"f8",
          3108 => x"c2",
          3109 => x"ec",
          3110 => x"98",
          3111 => x"53",
          3112 => x"51",
          3113 => x"82",
          3114 => x"81",
          3115 => x"73",
          3116 => x"38",
          3117 => x"81",
          3118 => x"54",
          3119 => x"ff",
          3120 => x"54",
          3121 => x"ec",
          3122 => x"0d",
          3123 => x"0d",
          3124 => x"b2",
          3125 => x"3d",
          3126 => x"5a",
          3127 => x"3d",
          3128 => x"c4",
          3129 => x"c0",
          3130 => x"73",
          3131 => x"73",
          3132 => x"33",
          3133 => x"83",
          3134 => x"76",
          3135 => x"bb",
          3136 => x"76",
          3137 => x"73",
          3138 => x"ac",
          3139 => x"97",
          3140 => x"85",
          3141 => x"85",
          3142 => x"85",
          3143 => x"2e",
          3144 => x"93",
          3145 => x"82",
          3146 => x"51",
          3147 => x"3f",
          3148 => x"08",
          3149 => x"38",
          3150 => x"51",
          3151 => x"80",
          3152 => x"85",
          3153 => x"82",
          3154 => x"53",
          3155 => x"90",
          3156 => x"54",
          3157 => x"3f",
          3158 => x"08",
          3159 => x"ec",
          3160 => x"09",
          3161 => x"d0",
          3162 => x"ec",
          3163 => x"b0",
          3164 => x"85",
          3165 => x"80",
          3166 => x"ec",
          3167 => x"38",
          3168 => x"08",
          3169 => x"17",
          3170 => x"74",
          3171 => x"74",
          3172 => x"52",
          3173 => x"c5",
          3174 => x"70",
          3175 => x"5c",
          3176 => x"27",
          3177 => x"5b",
          3178 => x"09",
          3179 => x"97",
          3180 => x"75",
          3181 => x"34",
          3182 => x"82",
          3183 => x"80",
          3184 => x"f9",
          3185 => x"3d",
          3186 => x"3f",
          3187 => x"08",
          3188 => x"98",
          3189 => x"78",
          3190 => x"38",
          3191 => x"06",
          3192 => x"33",
          3193 => x"70",
          3194 => x"9d",
          3195 => x"98",
          3196 => x"2c",
          3197 => x"05",
          3198 => x"81",
          3199 => x"08",
          3200 => x"51",
          3201 => x"59",
          3202 => x"5d",
          3203 => x"73",
          3204 => x"e3",
          3205 => x"27",
          3206 => x"15",
          3207 => x"70",
          3208 => x"56",
          3209 => x"24",
          3210 => x"76",
          3211 => x"77",
          3212 => x"3f",
          3213 => x"08",
          3214 => x"54",
          3215 => x"da",
          3216 => x"9d",
          3217 => x"56",
          3218 => x"15",
          3219 => x"70",
          3220 => x"81",
          3221 => x"51",
          3222 => x"95",
          3223 => x"76",
          3224 => x"77",
          3225 => x"3f",
          3226 => x"08",
          3227 => x"54",
          3228 => x"d6",
          3229 => x"75",
          3230 => x"ca",
          3231 => x"54",
          3232 => x"84",
          3233 => x"2b",
          3234 => x"82",
          3235 => x"70",
          3236 => x"98",
          3237 => x"71",
          3238 => x"81",
          3239 => x"33",
          3240 => x"51",
          3241 => x"54",
          3242 => x"09",
          3243 => x"99",
          3244 => x"fc",
          3245 => x"0c",
          3246 => x"9d",
          3247 => x"0b",
          3248 => x"34",
          3249 => x"82",
          3250 => x"75",
          3251 => x"34",
          3252 => x"34",
          3253 => x"7e",
          3254 => x"26",
          3255 => x"73",
          3256 => x"81",
          3257 => x"08",
          3258 => x"8c",
          3259 => x"7e",
          3260 => x"38",
          3261 => x"33",
          3262 => x"27",
          3263 => x"98",
          3264 => x"2c",
          3265 => x"75",
          3266 => x"74",
          3267 => x"33",
          3268 => x"ff",
          3269 => x"2b",
          3270 => x"82",
          3271 => x"53",
          3272 => x"74",
          3273 => x"38",
          3274 => x"33",
          3275 => x"54",
          3276 => x"8c",
          3277 => x"54",
          3278 => x"74",
          3279 => x"88",
          3280 => x"7e",
          3281 => x"81",
          3282 => x"82",
          3283 => x"82",
          3284 => x"ff",
          3285 => x"2b",
          3286 => x"82",
          3287 => x"59",
          3288 => x"74",
          3289 => x"38",
          3290 => x"33",
          3291 => x"a1",
          3292 => x"70",
          3293 => x"98",
          3294 => x"88",
          3295 => x"56",
          3296 => x"24",
          3297 => x"9d",
          3298 => x"98",
          3299 => x"2c",
          3300 => x"33",
          3301 => x"54",
          3302 => x"fc",
          3303 => x"51",
          3304 => x"81",
          3305 => x"2b",
          3306 => x"82",
          3307 => x"5a",
          3308 => x"76",
          3309 => x"38",
          3310 => x"83",
          3311 => x"0b",
          3312 => x"82",
          3313 => x"80",
          3314 => x"d8",
          3315 => x"3f",
          3316 => x"82",
          3317 => x"70",
          3318 => x"55",
          3319 => x"2e",
          3320 => x"82",
          3321 => x"ff",
          3322 => x"82",
          3323 => x"ff",
          3324 => x"82",
          3325 => x"88",
          3326 => x"3f",
          3327 => x"33",
          3328 => x"70",
          3329 => x"9d",
          3330 => x"51",
          3331 => x"74",
          3332 => x"74",
          3333 => x"14",
          3334 => x"73",
          3335 => x"f1",
          3336 => x"70",
          3337 => x"98",
          3338 => x"88",
          3339 => x"56",
          3340 => x"24",
          3341 => x"51",
          3342 => x"82",
          3343 => x"70",
          3344 => x"98",
          3345 => x"88",
          3346 => x"56",
          3347 => x"24",
          3348 => x"88",
          3349 => x"3f",
          3350 => x"98",
          3351 => x"2c",
          3352 => x"33",
          3353 => x"54",
          3354 => x"e7",
          3355 => x"39",
          3356 => x"33",
          3357 => x"80",
          3358 => x"51",
          3359 => x"82",
          3360 => x"79",
          3361 => x"3f",
          3362 => x"08",
          3363 => x"54",
          3364 => x"82",
          3365 => x"54",
          3366 => x"8f",
          3367 => x"73",
          3368 => x"f2",
          3369 => x"39",
          3370 => x"80",
          3371 => x"8c",
          3372 => x"82",
          3373 => x"79",
          3374 => x"0c",
          3375 => x"04",
          3376 => x"33",
          3377 => x"2e",
          3378 => x"88",
          3379 => x"3f",
          3380 => x"33",
          3381 => x"73",
          3382 => x"34",
          3383 => x"06",
          3384 => x"82",
          3385 => x"82",
          3386 => x"55",
          3387 => x"2e",
          3388 => x"ff",
          3389 => x"82",
          3390 => x"74",
          3391 => x"98",
          3392 => x"ff",
          3393 => x"55",
          3394 => x"a4",
          3395 => x"54",
          3396 => x"74",
          3397 => x"51",
          3398 => x"81",
          3399 => x"2b",
          3400 => x"82",
          3401 => x"59",
          3402 => x"75",
          3403 => x"38",
          3404 => x"dd",
          3405 => x"8c",
          3406 => x"2b",
          3407 => x"82",
          3408 => x"57",
          3409 => x"74",
          3410 => x"fa",
          3411 => x"e3",
          3412 => x"15",
          3413 => x"70",
          3414 => x"9d",
          3415 => x"51",
          3416 => x"75",
          3417 => x"f8",
          3418 => x"9d",
          3419 => x"81",
          3420 => x"9d",
          3421 => x"56",
          3422 => x"27",
          3423 => x"81",
          3424 => x"82",
          3425 => x"74",
          3426 => x"52",
          3427 => x"3f",
          3428 => x"33",
          3429 => x"06",
          3430 => x"33",
          3431 => x"75",
          3432 => x"38",
          3433 => x"82",
          3434 => x"80",
          3435 => x"d8",
          3436 => x"3f",
          3437 => x"9d",
          3438 => x"0b",
          3439 => x"34",
          3440 => x"7a",
          3441 => x"85",
          3442 => x"74",
          3443 => x"38",
          3444 => x"a7",
          3445 => x"85",
          3446 => x"9d",
          3447 => x"85",
          3448 => x"ff",
          3449 => x"53",
          3450 => x"51",
          3451 => x"3f",
          3452 => x"c0",
          3453 => x"2b",
          3454 => x"11",
          3455 => x"57",
          3456 => x"80",
          3457 => x"74",
          3458 => x"b0",
          3459 => x"ec",
          3460 => x"88",
          3461 => x"ec",
          3462 => x"06",
          3463 => x"74",
          3464 => x"ff",
          3465 => x"ff",
          3466 => x"f9",
          3467 => x"55",
          3468 => x"f7",
          3469 => x"51",
          3470 => x"3f",
          3471 => x"93",
          3472 => x"06",
          3473 => x"84",
          3474 => x"74",
          3475 => x"38",
          3476 => x"a6",
          3477 => x"85",
          3478 => x"9d",
          3479 => x"85",
          3480 => x"ff",
          3481 => x"53",
          3482 => x"51",
          3483 => x"3f",
          3484 => x"7a",
          3485 => x"84",
          3486 => x"56",
          3487 => x"2e",
          3488 => x"51",
          3489 => x"3f",
          3490 => x"08",
          3491 => x"34",
          3492 => x"08",
          3493 => x"81",
          3494 => x"52",
          3495 => x"a7",
          3496 => x"1b",
          3497 => x"ff",
          3498 => x"39",
          3499 => x"88",
          3500 => x"34",
          3501 => x"53",
          3502 => x"33",
          3503 => x"ed",
          3504 => x"82",
          3505 => x"8c",
          3506 => x"ff",
          3507 => x"88",
          3508 => x"54",
          3509 => x"f5",
          3510 => x"14",
          3511 => x"9d",
          3512 => x"1a",
          3513 => x"54",
          3514 => x"f5",
          3515 => x"9d",
          3516 => x"73",
          3517 => x"ce",
          3518 => x"e0",
          3519 => x"9d",
          3520 => x"05",
          3521 => x"9d",
          3522 => x"ba",
          3523 => x"0d",
          3524 => x"0b",
          3525 => x"0c",
          3526 => x"82",
          3527 => x"90",
          3528 => x"52",
          3529 => x"51",
          3530 => x"3f",
          3531 => x"08",
          3532 => x"77",
          3533 => x"57",
          3534 => x"34",
          3535 => x"08",
          3536 => x"15",
          3537 => x"15",
          3538 => x"e4",
          3539 => x"86",
          3540 => x"87",
          3541 => x"85",
          3542 => x"85",
          3543 => x"05",
          3544 => x"07",
          3545 => x"ff",
          3546 => x"2a",
          3547 => x"56",
          3548 => x"34",
          3549 => x"34",
          3550 => x"22",
          3551 => x"82",
          3552 => x"11",
          3553 => x"55",
          3554 => x"15",
          3555 => x"15",
          3556 => x"0d",
          3557 => x"0d",
          3558 => x"51",
          3559 => x"8f",
          3560 => x"83",
          3561 => x"70",
          3562 => x"06",
          3563 => x"70",
          3564 => x"0c",
          3565 => x"04",
          3566 => x"02",
          3567 => x"02",
          3568 => x"05",
          3569 => x"82",
          3570 => x"71",
          3571 => x"11",
          3572 => x"73",
          3573 => x"81",
          3574 => x"88",
          3575 => x"a4",
          3576 => x"22",
          3577 => x"ff",
          3578 => x"88",
          3579 => x"52",
          3580 => x"5b",
          3581 => x"55",
          3582 => x"70",
          3583 => x"82",
          3584 => x"14",
          3585 => x"52",
          3586 => x"15",
          3587 => x"15",
          3588 => x"e4",
          3589 => x"70",
          3590 => x"33",
          3591 => x"07",
          3592 => x"8f",
          3593 => x"51",
          3594 => x"71",
          3595 => x"ff",
          3596 => x"88",
          3597 => x"51",
          3598 => x"34",
          3599 => x"06",
          3600 => x"12",
          3601 => x"e4",
          3602 => x"71",
          3603 => x"81",
          3604 => x"3d",
          3605 => x"3d",
          3606 => x"e4",
          3607 => x"05",
          3608 => x"70",
          3609 => x"11",
          3610 => x"87",
          3611 => x"8b",
          3612 => x"2b",
          3613 => x"59",
          3614 => x"72",
          3615 => x"33",
          3616 => x"71",
          3617 => x"70",
          3618 => x"56",
          3619 => x"84",
          3620 => x"85",
          3621 => x"85",
          3622 => x"14",
          3623 => x"85",
          3624 => x"8b",
          3625 => x"2b",
          3626 => x"57",
          3627 => x"86",
          3628 => x"13",
          3629 => x"2b",
          3630 => x"2a",
          3631 => x"52",
          3632 => x"34",
          3633 => x"34",
          3634 => x"08",
          3635 => x"81",
          3636 => x"88",
          3637 => x"81",
          3638 => x"70",
          3639 => x"51",
          3640 => x"71",
          3641 => x"81",
          3642 => x"3d",
          3643 => x"3d",
          3644 => x"05",
          3645 => x"e4",
          3646 => x"2b",
          3647 => x"33",
          3648 => x"71",
          3649 => x"70",
          3650 => x"59",
          3651 => x"73",
          3652 => x"81",
          3653 => x"98",
          3654 => x"2b",
          3655 => x"55",
          3656 => x"80",
          3657 => x"38",
          3658 => x"aa",
          3659 => x"e4",
          3660 => x"70",
          3661 => x"33",
          3662 => x"71",
          3663 => x"74",
          3664 => x"81",
          3665 => x"88",
          3666 => x"83",
          3667 => x"f8",
          3668 => x"5d",
          3669 => x"5a",
          3670 => x"75",
          3671 => x"52",
          3672 => x"34",
          3673 => x"34",
          3674 => x"08",
          3675 => x"33",
          3676 => x"71",
          3677 => x"83",
          3678 => x"59",
          3679 => x"05",
          3680 => x"12",
          3681 => x"2b",
          3682 => x"ff",
          3683 => x"88",
          3684 => x"52",
          3685 => x"74",
          3686 => x"15",
          3687 => x"0d",
          3688 => x"0d",
          3689 => x"08",
          3690 => x"9e",
          3691 => x"83",
          3692 => x"82",
          3693 => x"12",
          3694 => x"2b",
          3695 => x"07",
          3696 => x"52",
          3697 => x"05",
          3698 => x"13",
          3699 => x"2b",
          3700 => x"05",
          3701 => x"71",
          3702 => x"2a",
          3703 => x"53",
          3704 => x"34",
          3705 => x"34",
          3706 => x"08",
          3707 => x"33",
          3708 => x"71",
          3709 => x"83",
          3710 => x"59",
          3711 => x"05",
          3712 => x"83",
          3713 => x"88",
          3714 => x"88",
          3715 => x"56",
          3716 => x"13",
          3717 => x"13",
          3718 => x"e4",
          3719 => x"11",
          3720 => x"33",
          3721 => x"07",
          3722 => x"0c",
          3723 => x"3d",
          3724 => x"3d",
          3725 => x"85",
          3726 => x"83",
          3727 => x"ff",
          3728 => x"53",
          3729 => x"a6",
          3730 => x"e4",
          3731 => x"2b",
          3732 => x"11",
          3733 => x"33",
          3734 => x"71",
          3735 => x"75",
          3736 => x"81",
          3737 => x"98",
          3738 => x"2b",
          3739 => x"40",
          3740 => x"58",
          3741 => x"72",
          3742 => x"38",
          3743 => x"52",
          3744 => x"9d",
          3745 => x"39",
          3746 => x"85",
          3747 => x"8b",
          3748 => x"2b",
          3749 => x"79",
          3750 => x"51",
          3751 => x"76",
          3752 => x"75",
          3753 => x"56",
          3754 => x"34",
          3755 => x"08",
          3756 => x"12",
          3757 => x"33",
          3758 => x"07",
          3759 => x"54",
          3760 => x"53",
          3761 => x"34",
          3762 => x"34",
          3763 => x"08",
          3764 => x"0b",
          3765 => x"80",
          3766 => x"34",
          3767 => x"08",
          3768 => x"14",
          3769 => x"14",
          3770 => x"e4",
          3771 => x"33",
          3772 => x"71",
          3773 => x"70",
          3774 => x"07",
          3775 => x"53",
          3776 => x"54",
          3777 => x"72",
          3778 => x"8b",
          3779 => x"ff",
          3780 => x"52",
          3781 => x"08",
          3782 => x"f1",
          3783 => x"2e",
          3784 => x"51",
          3785 => x"83",
          3786 => x"f5",
          3787 => x"7e",
          3788 => x"e1",
          3789 => x"ec",
          3790 => x"ff",
          3791 => x"e4",
          3792 => x"33",
          3793 => x"71",
          3794 => x"70",
          3795 => x"58",
          3796 => x"ff",
          3797 => x"2e",
          3798 => x"75",
          3799 => x"05",
          3800 => x"12",
          3801 => x"2b",
          3802 => x"ff",
          3803 => x"31",
          3804 => x"ff",
          3805 => x"27",
          3806 => x"56",
          3807 => x"79",
          3808 => x"73",
          3809 => x"38",
          3810 => x"5b",
          3811 => x"85",
          3812 => x"88",
          3813 => x"54",
          3814 => x"78",
          3815 => x"2e",
          3816 => x"79",
          3817 => x"76",
          3818 => x"85",
          3819 => x"70",
          3820 => x"33",
          3821 => x"07",
          3822 => x"ff",
          3823 => x"5a",
          3824 => x"73",
          3825 => x"38",
          3826 => x"54",
          3827 => x"81",
          3828 => x"54",
          3829 => x"81",
          3830 => x"7a",
          3831 => x"06",
          3832 => x"51",
          3833 => x"81",
          3834 => x"80",
          3835 => x"52",
          3836 => x"c4",
          3837 => x"e4",
          3838 => x"86",
          3839 => x"12",
          3840 => x"2b",
          3841 => x"07",
          3842 => x"55",
          3843 => x"17",
          3844 => x"ff",
          3845 => x"2a",
          3846 => x"54",
          3847 => x"34",
          3848 => x"06",
          3849 => x"15",
          3850 => x"e4",
          3851 => x"2b",
          3852 => x"1e",
          3853 => x"87",
          3854 => x"88",
          3855 => x"88",
          3856 => x"5e",
          3857 => x"54",
          3858 => x"34",
          3859 => x"34",
          3860 => x"08",
          3861 => x"11",
          3862 => x"33",
          3863 => x"71",
          3864 => x"53",
          3865 => x"74",
          3866 => x"86",
          3867 => x"87",
          3868 => x"85",
          3869 => x"16",
          3870 => x"11",
          3871 => x"33",
          3872 => x"07",
          3873 => x"53",
          3874 => x"56",
          3875 => x"16",
          3876 => x"16",
          3877 => x"e4",
          3878 => x"05",
          3879 => x"85",
          3880 => x"3d",
          3881 => x"3d",
          3882 => x"82",
          3883 => x"84",
          3884 => x"3f",
          3885 => x"80",
          3886 => x"71",
          3887 => x"3f",
          3888 => x"08",
          3889 => x"85",
          3890 => x"3d",
          3891 => x"3d",
          3892 => x"05",
          3893 => x"52",
          3894 => x"87",
          3895 => x"e8",
          3896 => x"71",
          3897 => x"0c",
          3898 => x"04",
          3899 => x"02",
          3900 => x"02",
          3901 => x"05",
          3902 => x"83",
          3903 => x"26",
          3904 => x"72",
          3905 => x"c0",
          3906 => x"53",
          3907 => x"74",
          3908 => x"38",
          3909 => x"73",
          3910 => x"c0",
          3911 => x"51",
          3912 => x"85",
          3913 => x"98",
          3914 => x"52",
          3915 => x"82",
          3916 => x"70",
          3917 => x"38",
          3918 => x"8c",
          3919 => x"ec",
          3920 => x"fc",
          3921 => x"52",
          3922 => x"87",
          3923 => x"08",
          3924 => x"2e",
          3925 => x"82",
          3926 => x"34",
          3927 => x"13",
          3928 => x"82",
          3929 => x"86",
          3930 => x"f3",
          3931 => x"62",
          3932 => x"05",
          3933 => x"57",
          3934 => x"83",
          3935 => x"fe",
          3936 => x"85",
          3937 => x"06",
          3938 => x"71",
          3939 => x"71",
          3940 => x"2b",
          3941 => x"80",
          3942 => x"92",
          3943 => x"c0",
          3944 => x"41",
          3945 => x"5a",
          3946 => x"87",
          3947 => x"0c",
          3948 => x"84",
          3949 => x"08",
          3950 => x"70",
          3951 => x"53",
          3952 => x"2e",
          3953 => x"08",
          3954 => x"70",
          3955 => x"34",
          3956 => x"80",
          3957 => x"53",
          3958 => x"2e",
          3959 => x"53",
          3960 => x"26",
          3961 => x"80",
          3962 => x"87",
          3963 => x"08",
          3964 => x"38",
          3965 => x"8c",
          3966 => x"80",
          3967 => x"78",
          3968 => x"99",
          3969 => x"0c",
          3970 => x"8c",
          3971 => x"08",
          3972 => x"51",
          3973 => x"38",
          3974 => x"8d",
          3975 => x"17",
          3976 => x"81",
          3977 => x"53",
          3978 => x"2e",
          3979 => x"fc",
          3980 => x"52",
          3981 => x"7d",
          3982 => x"ed",
          3983 => x"80",
          3984 => x"71",
          3985 => x"38",
          3986 => x"53",
          3987 => x"ec",
          3988 => x"0d",
          3989 => x"0d",
          3990 => x"02",
          3991 => x"05",
          3992 => x"58",
          3993 => x"80",
          3994 => x"fc",
          3995 => x"85",
          3996 => x"06",
          3997 => x"71",
          3998 => x"81",
          3999 => x"38",
          4000 => x"2b",
          4001 => x"80",
          4002 => x"92",
          4003 => x"c0",
          4004 => x"40",
          4005 => x"5a",
          4006 => x"c0",
          4007 => x"76",
          4008 => x"76",
          4009 => x"75",
          4010 => x"2a",
          4011 => x"51",
          4012 => x"80",
          4013 => x"7a",
          4014 => x"5c",
          4015 => x"81",
          4016 => x"81",
          4017 => x"06",
          4018 => x"80",
          4019 => x"87",
          4020 => x"08",
          4021 => x"38",
          4022 => x"8c",
          4023 => x"80",
          4024 => x"77",
          4025 => x"99",
          4026 => x"0c",
          4027 => x"8c",
          4028 => x"08",
          4029 => x"51",
          4030 => x"38",
          4031 => x"8d",
          4032 => x"70",
          4033 => x"84",
          4034 => x"5b",
          4035 => x"2e",
          4036 => x"fc",
          4037 => x"52",
          4038 => x"7d",
          4039 => x"f8",
          4040 => x"80",
          4041 => x"71",
          4042 => x"38",
          4043 => x"53",
          4044 => x"ec",
          4045 => x"0d",
          4046 => x"0d",
          4047 => x"05",
          4048 => x"02",
          4049 => x"05",
          4050 => x"54",
          4051 => x"fe",
          4052 => x"ec",
          4053 => x"53",
          4054 => x"80",
          4055 => x"0b",
          4056 => x"8c",
          4057 => x"71",
          4058 => x"dc",
          4059 => x"24",
          4060 => x"84",
          4061 => x"92",
          4062 => x"54",
          4063 => x"8d",
          4064 => x"39",
          4065 => x"80",
          4066 => x"cb",
          4067 => x"70",
          4068 => x"81",
          4069 => x"52",
          4070 => x"8a",
          4071 => x"98",
          4072 => x"71",
          4073 => x"c0",
          4074 => x"52",
          4075 => x"81",
          4076 => x"c0",
          4077 => x"53",
          4078 => x"82",
          4079 => x"71",
          4080 => x"39",
          4081 => x"39",
          4082 => x"77",
          4083 => x"81",
          4084 => x"72",
          4085 => x"84",
          4086 => x"73",
          4087 => x"0c",
          4088 => x"04",
          4089 => x"74",
          4090 => x"71",
          4091 => x"2b",
          4092 => x"ec",
          4093 => x"84",
          4094 => x"fd",
          4095 => x"83",
          4096 => x"12",
          4097 => x"2b",
          4098 => x"07",
          4099 => x"70",
          4100 => x"2b",
          4101 => x"07",
          4102 => x"0c",
          4103 => x"56",
          4104 => x"3d",
          4105 => x"3d",
          4106 => x"84",
          4107 => x"22",
          4108 => x"72",
          4109 => x"54",
          4110 => x"2a",
          4111 => x"34",
          4112 => x"04",
          4113 => x"73",
          4114 => x"70",
          4115 => x"05",
          4116 => x"88",
          4117 => x"72",
          4118 => x"54",
          4119 => x"2a",
          4120 => x"70",
          4121 => x"34",
          4122 => x"51",
          4123 => x"83",
          4124 => x"fe",
          4125 => x"75",
          4126 => x"51",
          4127 => x"92",
          4128 => x"81",
          4129 => x"73",
          4130 => x"55",
          4131 => x"51",
          4132 => x"3d",
          4133 => x"3d",
          4134 => x"76",
          4135 => x"72",
          4136 => x"05",
          4137 => x"11",
          4138 => x"38",
          4139 => x"04",
          4140 => x"78",
          4141 => x"56",
          4142 => x"81",
          4143 => x"74",
          4144 => x"56",
          4145 => x"31",
          4146 => x"52",
          4147 => x"80",
          4148 => x"71",
          4149 => x"38",
          4150 => x"ec",
          4151 => x"0d",
          4152 => x"0d",
          4153 => x"51",
          4154 => x"73",
          4155 => x"81",
          4156 => x"33",
          4157 => x"38",
          4158 => x"85",
          4159 => x"3d",
          4160 => x"0b",
          4161 => x"0c",
          4162 => x"82",
          4163 => x"04",
          4164 => x"7b",
          4165 => x"83",
          4166 => x"5a",
          4167 => x"80",
          4168 => x"54",
          4169 => x"53",
          4170 => x"53",
          4171 => x"52",
          4172 => x"3f",
          4173 => x"08",
          4174 => x"81",
          4175 => x"82",
          4176 => x"83",
          4177 => x"16",
          4178 => x"18",
          4179 => x"18",
          4180 => x"58",
          4181 => x"9f",
          4182 => x"33",
          4183 => x"2e",
          4184 => x"93",
          4185 => x"76",
          4186 => x"52",
          4187 => x"51",
          4188 => x"83",
          4189 => x"79",
          4190 => x"0c",
          4191 => x"04",
          4192 => x"78",
          4193 => x"80",
          4194 => x"17",
          4195 => x"38",
          4196 => x"fc",
          4197 => x"ec",
          4198 => x"85",
          4199 => x"38",
          4200 => x"53",
          4201 => x"81",
          4202 => x"f7",
          4203 => x"85",
          4204 => x"2e",
          4205 => x"55",
          4206 => x"b0",
          4207 => x"82",
          4208 => x"88",
          4209 => x"f8",
          4210 => x"70",
          4211 => x"c0",
          4212 => x"ec",
          4213 => x"85",
          4214 => x"91",
          4215 => x"55",
          4216 => x"09",
          4217 => x"f0",
          4218 => x"33",
          4219 => x"2e",
          4220 => x"80",
          4221 => x"80",
          4222 => x"ec",
          4223 => x"17",
          4224 => x"fd",
          4225 => x"d4",
          4226 => x"b2",
          4227 => x"96",
          4228 => x"85",
          4229 => x"75",
          4230 => x"3f",
          4231 => x"e4",
          4232 => x"98",
          4233 => x"9c",
          4234 => x"08",
          4235 => x"17",
          4236 => x"3f",
          4237 => x"52",
          4238 => x"51",
          4239 => x"a0",
          4240 => x"05",
          4241 => x"0c",
          4242 => x"75",
          4243 => x"33",
          4244 => x"3f",
          4245 => x"34",
          4246 => x"52",
          4247 => x"51",
          4248 => x"82",
          4249 => x"80",
          4250 => x"81",
          4251 => x"85",
          4252 => x"3d",
          4253 => x"3d",
          4254 => x"1a",
          4255 => x"fe",
          4256 => x"55",
          4257 => x"73",
          4258 => x"8a",
          4259 => x"53",
          4260 => x"f9",
          4261 => x"08",
          4262 => x"08",
          4263 => x"82",
          4264 => x"87",
          4265 => x"f9",
          4266 => x"7a",
          4267 => x"54",
          4268 => x"27",
          4269 => x"76",
          4270 => x"27",
          4271 => x"ff",
          4272 => x"58",
          4273 => x"80",
          4274 => x"82",
          4275 => x"72",
          4276 => x"38",
          4277 => x"72",
          4278 => x"8e",
          4279 => x"39",
          4280 => x"17",
          4281 => x"a4",
          4282 => x"53",
          4283 => x"fd",
          4284 => x"85",
          4285 => x"9f",
          4286 => x"ff",
          4287 => x"11",
          4288 => x"70",
          4289 => x"18",
          4290 => x"76",
          4291 => x"53",
          4292 => x"82",
          4293 => x"80",
          4294 => x"83",
          4295 => x"b4",
          4296 => x"88",
          4297 => x"79",
          4298 => x"84",
          4299 => x"58",
          4300 => x"80",
          4301 => x"9f",
          4302 => x"80",
          4303 => x"88",
          4304 => x"08",
          4305 => x"51",
          4306 => x"82",
          4307 => x"80",
          4308 => x"10",
          4309 => x"74",
          4310 => x"51",
          4311 => x"82",
          4312 => x"83",
          4313 => x"58",
          4314 => x"87",
          4315 => x"08",
          4316 => x"51",
          4317 => x"82",
          4318 => x"9b",
          4319 => x"2b",
          4320 => x"74",
          4321 => x"51",
          4322 => x"82",
          4323 => x"f0",
          4324 => x"83",
          4325 => x"77",
          4326 => x"0c",
          4327 => x"04",
          4328 => x"7a",
          4329 => x"58",
          4330 => x"81",
          4331 => x"9e",
          4332 => x"17",
          4333 => x"96",
          4334 => x"53",
          4335 => x"81",
          4336 => x"79",
          4337 => x"72",
          4338 => x"38",
          4339 => x"72",
          4340 => x"b8",
          4341 => x"39",
          4342 => x"17",
          4343 => x"a4",
          4344 => x"53",
          4345 => x"fb",
          4346 => x"85",
          4347 => x"82",
          4348 => x"81",
          4349 => x"83",
          4350 => x"b4",
          4351 => x"78",
          4352 => x"56",
          4353 => x"76",
          4354 => x"38",
          4355 => x"9f",
          4356 => x"33",
          4357 => x"07",
          4358 => x"74",
          4359 => x"83",
          4360 => x"89",
          4361 => x"08",
          4362 => x"51",
          4363 => x"82",
          4364 => x"59",
          4365 => x"08",
          4366 => x"74",
          4367 => x"16",
          4368 => x"84",
          4369 => x"76",
          4370 => x"88",
          4371 => x"81",
          4372 => x"8f",
          4373 => x"53",
          4374 => x"80",
          4375 => x"88",
          4376 => x"08",
          4377 => x"51",
          4378 => x"82",
          4379 => x"59",
          4380 => x"08",
          4381 => x"77",
          4382 => x"06",
          4383 => x"83",
          4384 => x"05",
          4385 => x"f7",
          4386 => x"39",
          4387 => x"a4",
          4388 => x"52",
          4389 => x"e8",
          4390 => x"ec",
          4391 => x"85",
          4392 => x"38",
          4393 => x"06",
          4394 => x"83",
          4395 => x"18",
          4396 => x"54",
          4397 => x"f6",
          4398 => x"85",
          4399 => x"0a",
          4400 => x"52",
          4401 => x"fc",
          4402 => x"83",
          4403 => x"82",
          4404 => x"8a",
          4405 => x"f8",
          4406 => x"7c",
          4407 => x"59",
          4408 => x"81",
          4409 => x"38",
          4410 => x"08",
          4411 => x"73",
          4412 => x"38",
          4413 => x"52",
          4414 => x"a4",
          4415 => x"ec",
          4416 => x"85",
          4417 => x"f2",
          4418 => x"82",
          4419 => x"39",
          4420 => x"e6",
          4421 => x"ec",
          4422 => x"de",
          4423 => x"78",
          4424 => x"3f",
          4425 => x"08",
          4426 => x"ec",
          4427 => x"80",
          4428 => x"85",
          4429 => x"2e",
          4430 => x"85",
          4431 => x"2e",
          4432 => x"53",
          4433 => x"51",
          4434 => x"82",
          4435 => x"c5",
          4436 => x"08",
          4437 => x"18",
          4438 => x"57",
          4439 => x"90",
          4440 => x"90",
          4441 => x"16",
          4442 => x"54",
          4443 => x"34",
          4444 => x"78",
          4445 => x"38",
          4446 => x"82",
          4447 => x"8a",
          4448 => x"f6",
          4449 => x"7e",
          4450 => x"5b",
          4451 => x"38",
          4452 => x"58",
          4453 => x"88",
          4454 => x"08",
          4455 => x"38",
          4456 => x"39",
          4457 => x"51",
          4458 => x"81",
          4459 => x"85",
          4460 => x"82",
          4461 => x"85",
          4462 => x"82",
          4463 => x"ff",
          4464 => x"38",
          4465 => x"82",
          4466 => x"26",
          4467 => x"79",
          4468 => x"08",
          4469 => x"73",
          4470 => x"bf",
          4471 => x"2e",
          4472 => x"80",
          4473 => x"1a",
          4474 => x"08",
          4475 => x"38",
          4476 => x"52",
          4477 => x"af",
          4478 => x"82",
          4479 => x"81",
          4480 => x"06",
          4481 => x"85",
          4482 => x"82",
          4483 => x"09",
          4484 => x"05",
          4485 => x"80",
          4486 => x"07",
          4487 => x"08",
          4488 => x"55",
          4489 => x"f3",
          4490 => x"ec",
          4491 => x"95",
          4492 => x"08",
          4493 => x"27",
          4494 => x"98",
          4495 => x"89",
          4496 => x"85",
          4497 => x"dd",
          4498 => x"81",
          4499 => x"17",
          4500 => x"89",
          4501 => x"75",
          4502 => x"b0",
          4503 => x"7a",
          4504 => x"3f",
          4505 => x"08",
          4506 => x"38",
          4507 => x"85",
          4508 => x"2e",
          4509 => x"86",
          4510 => x"ec",
          4511 => x"85",
          4512 => x"70",
          4513 => x"70",
          4514 => x"25",
          4515 => x"51",
          4516 => x"73",
          4517 => x"75",
          4518 => x"81",
          4519 => x"38",
          4520 => x"f7",
          4521 => x"75",
          4522 => x"f9",
          4523 => x"85",
          4524 => x"85",
          4525 => x"81",
          4526 => x"85",
          4527 => x"80",
          4528 => x"55",
          4529 => x"94",
          4530 => x"2e",
          4531 => x"53",
          4532 => x"51",
          4533 => x"82",
          4534 => x"55",
          4535 => x"75",
          4536 => x"98",
          4537 => x"05",
          4538 => x"56",
          4539 => x"26",
          4540 => x"15",
          4541 => x"84",
          4542 => x"07",
          4543 => x"18",
          4544 => x"ff",
          4545 => x"2e",
          4546 => x"39",
          4547 => x"39",
          4548 => x"08",
          4549 => x"81",
          4550 => x"74",
          4551 => x"0c",
          4552 => x"04",
          4553 => x"7a",
          4554 => x"f3",
          4555 => x"85",
          4556 => x"81",
          4557 => x"ec",
          4558 => x"38",
          4559 => x"51",
          4560 => x"82",
          4561 => x"82",
          4562 => x"b0",
          4563 => x"84",
          4564 => x"52",
          4565 => x"52",
          4566 => x"3f",
          4567 => x"39",
          4568 => x"8a",
          4569 => x"75",
          4570 => x"38",
          4571 => x"19",
          4572 => x"81",
          4573 => x"ed",
          4574 => x"85",
          4575 => x"2e",
          4576 => x"15",
          4577 => x"70",
          4578 => x"70",
          4579 => x"9f",
          4580 => x"56",
          4581 => x"85",
          4582 => x"3d",
          4583 => x"3d",
          4584 => x"71",
          4585 => x"57",
          4586 => x"0a",
          4587 => x"38",
          4588 => x"53",
          4589 => x"38",
          4590 => x"0c",
          4591 => x"54",
          4592 => x"75",
          4593 => x"73",
          4594 => x"a8",
          4595 => x"73",
          4596 => x"85",
          4597 => x"0b",
          4598 => x"5a",
          4599 => x"27",
          4600 => x"a8",
          4601 => x"18",
          4602 => x"39",
          4603 => x"70",
          4604 => x"58",
          4605 => x"b2",
          4606 => x"76",
          4607 => x"3f",
          4608 => x"08",
          4609 => x"ec",
          4610 => x"bd",
          4611 => x"82",
          4612 => x"27",
          4613 => x"16",
          4614 => x"ec",
          4615 => x"38",
          4616 => x"39",
          4617 => x"55",
          4618 => x"52",
          4619 => x"c6",
          4620 => x"ec",
          4621 => x"0c",
          4622 => x"0c",
          4623 => x"53",
          4624 => x"80",
          4625 => x"85",
          4626 => x"94",
          4627 => x"2a",
          4628 => x"0c",
          4629 => x"06",
          4630 => x"9c",
          4631 => x"58",
          4632 => x"ec",
          4633 => x"0d",
          4634 => x"0d",
          4635 => x"90",
          4636 => x"05",
          4637 => x"f0",
          4638 => x"27",
          4639 => x"0b",
          4640 => x"98",
          4641 => x"84",
          4642 => x"2e",
          4643 => x"76",
          4644 => x"58",
          4645 => x"38",
          4646 => x"15",
          4647 => x"08",
          4648 => x"38",
          4649 => x"88",
          4650 => x"53",
          4651 => x"81",
          4652 => x"c0",
          4653 => x"22",
          4654 => x"89",
          4655 => x"72",
          4656 => x"74",
          4657 => x"f3",
          4658 => x"85",
          4659 => x"82",
          4660 => x"82",
          4661 => x"27",
          4662 => x"81",
          4663 => x"ec",
          4664 => x"80",
          4665 => x"16",
          4666 => x"ec",
          4667 => x"ca",
          4668 => x"38",
          4669 => x"0c",
          4670 => x"dd",
          4671 => x"08",
          4672 => x"f8",
          4673 => x"85",
          4674 => x"87",
          4675 => x"ec",
          4676 => x"80",
          4677 => x"55",
          4678 => x"08",
          4679 => x"38",
          4680 => x"85",
          4681 => x"2e",
          4682 => x"85",
          4683 => x"75",
          4684 => x"3f",
          4685 => x"08",
          4686 => x"94",
          4687 => x"52",
          4688 => x"b2",
          4689 => x"ec",
          4690 => x"0c",
          4691 => x"0c",
          4692 => x"05",
          4693 => x"80",
          4694 => x"85",
          4695 => x"3d",
          4696 => x"3d",
          4697 => x"71",
          4698 => x"57",
          4699 => x"51",
          4700 => x"82",
          4701 => x"54",
          4702 => x"08",
          4703 => x"82",
          4704 => x"56",
          4705 => x"52",
          4706 => x"f4",
          4707 => x"ec",
          4708 => x"85",
          4709 => x"d2",
          4710 => x"ec",
          4711 => x"08",
          4712 => x"54",
          4713 => x"e5",
          4714 => x"06",
          4715 => x"58",
          4716 => x"08",
          4717 => x"38",
          4718 => x"75",
          4719 => x"80",
          4720 => x"81",
          4721 => x"7a",
          4722 => x"06",
          4723 => x"39",
          4724 => x"08",
          4725 => x"76",
          4726 => x"3f",
          4727 => x"08",
          4728 => x"ec",
          4729 => x"ff",
          4730 => x"84",
          4731 => x"06",
          4732 => x"54",
          4733 => x"ec",
          4734 => x"0d",
          4735 => x"0d",
          4736 => x"52",
          4737 => x"3f",
          4738 => x"08",
          4739 => x"06",
          4740 => x"51",
          4741 => x"83",
          4742 => x"06",
          4743 => x"14",
          4744 => x"3f",
          4745 => x"08",
          4746 => x"07",
          4747 => x"85",
          4748 => x"3d",
          4749 => x"3d",
          4750 => x"70",
          4751 => x"06",
          4752 => x"53",
          4753 => x"de",
          4754 => x"33",
          4755 => x"83",
          4756 => x"06",
          4757 => x"90",
          4758 => x"15",
          4759 => x"3f",
          4760 => x"04",
          4761 => x"7b",
          4762 => x"84",
          4763 => x"58",
          4764 => x"80",
          4765 => x"38",
          4766 => x"52",
          4767 => x"80",
          4768 => x"ec",
          4769 => x"85",
          4770 => x"f5",
          4771 => x"08",
          4772 => x"53",
          4773 => x"84",
          4774 => x"39",
          4775 => x"70",
          4776 => x"81",
          4777 => x"51",
          4778 => x"16",
          4779 => x"ec",
          4780 => x"81",
          4781 => x"38",
          4782 => x"ae",
          4783 => x"81",
          4784 => x"54",
          4785 => x"2e",
          4786 => x"8f",
          4787 => x"82",
          4788 => x"76",
          4789 => x"54",
          4790 => x"09",
          4791 => x"38",
          4792 => x"7a",
          4793 => x"80",
          4794 => x"fa",
          4795 => x"85",
          4796 => x"82",
          4797 => x"89",
          4798 => x"08",
          4799 => x"86",
          4800 => x"98",
          4801 => x"82",
          4802 => x"8b",
          4803 => x"fb",
          4804 => x"70",
          4805 => x"81",
          4806 => x"fc",
          4807 => x"85",
          4808 => x"82",
          4809 => x"b4",
          4810 => x"08",
          4811 => x"ec",
          4812 => x"85",
          4813 => x"82",
          4814 => x"a0",
          4815 => x"82",
          4816 => x"52",
          4817 => x"51",
          4818 => x"8b",
          4819 => x"52",
          4820 => x"51",
          4821 => x"81",
          4822 => x"34",
          4823 => x"ec",
          4824 => x"0d",
          4825 => x"0d",
          4826 => x"98",
          4827 => x"70",
          4828 => x"ec",
          4829 => x"85",
          4830 => x"38",
          4831 => x"53",
          4832 => x"81",
          4833 => x"34",
          4834 => x"04",
          4835 => x"78",
          4836 => x"80",
          4837 => x"34",
          4838 => x"80",
          4839 => x"38",
          4840 => x"18",
          4841 => x"9c",
          4842 => x"70",
          4843 => x"56",
          4844 => x"a0",
          4845 => x"71",
          4846 => x"81",
          4847 => x"81",
          4848 => x"89",
          4849 => x"06",
          4850 => x"73",
          4851 => x"55",
          4852 => x"55",
          4853 => x"81",
          4854 => x"81",
          4855 => x"74",
          4856 => x"75",
          4857 => x"52",
          4858 => x"13",
          4859 => x"08",
          4860 => x"33",
          4861 => x"9c",
          4862 => x"11",
          4863 => x"fb",
          4864 => x"ec",
          4865 => x"96",
          4866 => x"d8",
          4867 => x"ec",
          4868 => x"23",
          4869 => x"e7",
          4870 => x"85",
          4871 => x"17",
          4872 => x"0d",
          4873 => x"0d",
          4874 => x"5e",
          4875 => x"70",
          4876 => x"55",
          4877 => x"83",
          4878 => x"73",
          4879 => x"91",
          4880 => x"2e",
          4881 => x"1d",
          4882 => x"0c",
          4883 => x"15",
          4884 => x"70",
          4885 => x"56",
          4886 => x"09",
          4887 => x"38",
          4888 => x"80",
          4889 => x"09",
          4890 => x"80",
          4891 => x"51",
          4892 => x"da",
          4893 => x"1c",
          4894 => x"33",
          4895 => x"9f",
          4896 => x"ff",
          4897 => x"1c",
          4898 => x"7a",
          4899 => x"3f",
          4900 => x"08",
          4901 => x"39",
          4902 => x"a0",
          4903 => x"5e",
          4904 => x"52",
          4905 => x"ee",
          4906 => x"59",
          4907 => x"33",
          4908 => x"ae",
          4909 => x"06",
          4910 => x"78",
          4911 => x"81",
          4912 => x"32",
          4913 => x"05",
          4914 => x"73",
          4915 => x"51",
          4916 => x"57",
          4917 => x"38",
          4918 => x"75",
          4919 => x"17",
          4920 => x"75",
          4921 => x"09",
          4922 => x"9f",
          4923 => x"54",
          4924 => x"2e",
          4925 => x"80",
          4926 => x"75",
          4927 => x"c7",
          4928 => x"7e",
          4929 => x"a0",
          4930 => x"c7",
          4931 => x"82",
          4932 => x"18",
          4933 => x"1a",
          4934 => x"a0",
          4935 => x"86",
          4936 => x"32",
          4937 => x"05",
          4938 => x"32",
          4939 => x"05",
          4940 => x"71",
          4941 => x"51",
          4942 => x"55",
          4943 => x"ae",
          4944 => x"81",
          4945 => x"78",
          4946 => x"51",
          4947 => x"af",
          4948 => x"06",
          4949 => x"55",
          4950 => x"32",
          4951 => x"05",
          4952 => x"77",
          4953 => x"54",
          4954 => x"81",
          4955 => x"ae",
          4956 => x"06",
          4957 => x"54",
          4958 => x"74",
          4959 => x"80",
          4960 => x"7b",
          4961 => x"09",
          4962 => x"ae",
          4963 => x"81",
          4964 => x"25",
          4965 => x"07",
          4966 => x"51",
          4967 => x"a7",
          4968 => x"8b",
          4969 => x"39",
          4970 => x"54",
          4971 => x"8c",
          4972 => x"ff",
          4973 => x"b4",
          4974 => x"54",
          4975 => x"c2",
          4976 => x"ec",
          4977 => x"b2",
          4978 => x"70",
          4979 => x"71",
          4980 => x"54",
          4981 => x"82",
          4982 => x"80",
          4983 => x"38",
          4984 => x"76",
          4985 => x"df",
          4986 => x"54",
          4987 => x"81",
          4988 => x"55",
          4989 => x"34",
          4990 => x"52",
          4991 => x"51",
          4992 => x"82",
          4993 => x"bf",
          4994 => x"16",
          4995 => x"26",
          4996 => x"16",
          4997 => x"06",
          4998 => x"17",
          4999 => x"34",
          5000 => x"fd",
          5001 => x"19",
          5002 => x"80",
          5003 => x"79",
          5004 => x"81",
          5005 => x"81",
          5006 => x"85",
          5007 => x"54",
          5008 => x"8f",
          5009 => x"86",
          5010 => x"39",
          5011 => x"f3",
          5012 => x"73",
          5013 => x"80",
          5014 => x"52",
          5015 => x"be",
          5016 => x"ec",
          5017 => x"85",
          5018 => x"d7",
          5019 => x"08",
          5020 => x"e6",
          5021 => x"85",
          5022 => x"82",
          5023 => x"80",
          5024 => x"1b",
          5025 => x"55",
          5026 => x"2e",
          5027 => x"8b",
          5028 => x"06",
          5029 => x"1c",
          5030 => x"33",
          5031 => x"70",
          5032 => x"55",
          5033 => x"38",
          5034 => x"52",
          5035 => x"80",
          5036 => x"ec",
          5037 => x"8b",
          5038 => x"7a",
          5039 => x"3f",
          5040 => x"75",
          5041 => x"57",
          5042 => x"2e",
          5043 => x"84",
          5044 => x"06",
          5045 => x"75",
          5046 => x"81",
          5047 => x"2a",
          5048 => x"73",
          5049 => x"38",
          5050 => x"54",
          5051 => x"fb",
          5052 => x"80",
          5053 => x"34",
          5054 => x"c1",
          5055 => x"06",
          5056 => x"38",
          5057 => x"39",
          5058 => x"70",
          5059 => x"54",
          5060 => x"86",
          5061 => x"84",
          5062 => x"06",
          5063 => x"73",
          5064 => x"38",
          5065 => x"83",
          5066 => x"b4",
          5067 => x"51",
          5068 => x"82",
          5069 => x"88",
          5070 => x"dc",
          5071 => x"85",
          5072 => x"3d",
          5073 => x"3d",
          5074 => x"ff",
          5075 => x"71",
          5076 => x"5c",
          5077 => x"80",
          5078 => x"38",
          5079 => x"05",
          5080 => x"a0",
          5081 => x"71",
          5082 => x"38",
          5083 => x"71",
          5084 => x"81",
          5085 => x"38",
          5086 => x"11",
          5087 => x"06",
          5088 => x"70",
          5089 => x"38",
          5090 => x"81",
          5091 => x"05",
          5092 => x"76",
          5093 => x"38",
          5094 => x"ff",
          5095 => x"77",
          5096 => x"57",
          5097 => x"05",
          5098 => x"70",
          5099 => x"33",
          5100 => x"53",
          5101 => x"99",
          5102 => x"e0",
          5103 => x"ff",
          5104 => x"ff",
          5105 => x"70",
          5106 => x"38",
          5107 => x"81",
          5108 => x"51",
          5109 => x"05",
          5110 => x"51",
          5111 => x"2e",
          5112 => x"85",
          5113 => x"bc",
          5114 => x"81",
          5115 => x"32",
          5116 => x"05",
          5117 => x"9f",
          5118 => x"2a",
          5119 => x"54",
          5120 => x"2e",
          5121 => x"15",
          5122 => x"55",
          5123 => x"ff",
          5124 => x"39",
          5125 => x"86",
          5126 => x"7c",
          5127 => x"51",
          5128 => x"9d",
          5129 => x"70",
          5130 => x"0c",
          5131 => x"04",
          5132 => x"78",
          5133 => x"83",
          5134 => x"0b",
          5135 => x"79",
          5136 => x"e2",
          5137 => x"55",
          5138 => x"08",
          5139 => x"84",
          5140 => x"df",
          5141 => x"85",
          5142 => x"ff",
          5143 => x"83",
          5144 => x"d4",
          5145 => x"81",
          5146 => x"38",
          5147 => x"17",
          5148 => x"74",
          5149 => x"09",
          5150 => x"38",
          5151 => x"81",
          5152 => x"09",
          5153 => x"80",
          5154 => x"51",
          5155 => x"8a",
          5156 => x"e8",
          5157 => x"06",
          5158 => x"53",
          5159 => x"52",
          5160 => x"51",
          5161 => x"82",
          5162 => x"55",
          5163 => x"08",
          5164 => x"38",
          5165 => x"fe",
          5166 => x"86",
          5167 => x"f0",
          5168 => x"ec",
          5169 => x"85",
          5170 => x"2e",
          5171 => x"55",
          5172 => x"ec",
          5173 => x"0d",
          5174 => x"0d",
          5175 => x"05",
          5176 => x"33",
          5177 => x"75",
          5178 => x"fc",
          5179 => x"85",
          5180 => x"8b",
          5181 => x"82",
          5182 => x"24",
          5183 => x"82",
          5184 => x"82",
          5185 => x"90",
          5186 => x"53",
          5187 => x"80",
          5188 => x"38",
          5189 => x"76",
          5190 => x"74",
          5191 => x"72",
          5192 => x"38",
          5193 => x"51",
          5194 => x"82",
          5195 => x"81",
          5196 => x"81",
          5197 => x"72",
          5198 => x"80",
          5199 => x"38",
          5200 => x"70",
          5201 => x"53",
          5202 => x"86",
          5203 => x"af",
          5204 => x"34",
          5205 => x"34",
          5206 => x"14",
          5207 => x"8c",
          5208 => x"ec",
          5209 => x"06",
          5210 => x"54",
          5211 => x"72",
          5212 => x"76",
          5213 => x"38",
          5214 => x"70",
          5215 => x"53",
          5216 => x"85",
          5217 => x"70",
          5218 => x"5c",
          5219 => x"82",
          5220 => x"81",
          5221 => x"76",
          5222 => x"81",
          5223 => x"38",
          5224 => x"56",
          5225 => x"83",
          5226 => x"70",
          5227 => x"80",
          5228 => x"83",
          5229 => x"dc",
          5230 => x"85",
          5231 => x"76",
          5232 => x"05",
          5233 => x"16",
          5234 => x"56",
          5235 => x"d7",
          5236 => x"8e",
          5237 => x"72",
          5238 => x"54",
          5239 => x"57",
          5240 => x"95",
          5241 => x"73",
          5242 => x"3f",
          5243 => x"08",
          5244 => x"57",
          5245 => x"89",
          5246 => x"56",
          5247 => x"d7",
          5248 => x"76",
          5249 => x"f9",
          5250 => x"76",
          5251 => x"f1",
          5252 => x"51",
          5253 => x"82",
          5254 => x"83",
          5255 => x"53",
          5256 => x"2e",
          5257 => x"84",
          5258 => x"ca",
          5259 => x"b4",
          5260 => x"ec",
          5261 => x"ff",
          5262 => x"8d",
          5263 => x"14",
          5264 => x"3f",
          5265 => x"08",
          5266 => x"15",
          5267 => x"14",
          5268 => x"34",
          5269 => x"33",
          5270 => x"81",
          5271 => x"54",
          5272 => x"72",
          5273 => x"99",
          5274 => x"ff",
          5275 => x"51",
          5276 => x"3f",
          5277 => x"08",
          5278 => x"33",
          5279 => x"8a",
          5280 => x"80",
          5281 => x"ff",
          5282 => x"53",
          5283 => x"86",
          5284 => x"83",
          5285 => x"c5",
          5286 => x"c8",
          5287 => x"ec",
          5288 => x"85",
          5289 => x"15",
          5290 => x"06",
          5291 => x"76",
          5292 => x"80",
          5293 => x"da",
          5294 => x"85",
          5295 => x"ff",
          5296 => x"74",
          5297 => x"d4",
          5298 => x"af",
          5299 => x"ec",
          5300 => x"c2",
          5301 => x"8c",
          5302 => x"ec",
          5303 => x"ff",
          5304 => x"56",
          5305 => x"83",
          5306 => x"14",
          5307 => x"71",
          5308 => x"5a",
          5309 => x"26",
          5310 => x"8a",
          5311 => x"74",
          5312 => x"fe",
          5313 => x"82",
          5314 => x"53",
          5315 => x"08",
          5316 => x"ed",
          5317 => x"ec",
          5318 => x"ff",
          5319 => x"83",
          5320 => x"72",
          5321 => x"26",
          5322 => x"57",
          5323 => x"26",
          5324 => x"57",
          5325 => x"56",
          5326 => x"82",
          5327 => x"13",
          5328 => x"0c",
          5329 => x"0c",
          5330 => x"a4",
          5331 => x"1e",
          5332 => x"54",
          5333 => x"2e",
          5334 => x"af",
          5335 => x"14",
          5336 => x"3f",
          5337 => x"08",
          5338 => x"06",
          5339 => x"72",
          5340 => x"7a",
          5341 => x"80",
          5342 => x"d8",
          5343 => x"85",
          5344 => x"15",
          5345 => x"2b",
          5346 => x"8d",
          5347 => x"2e",
          5348 => x"77",
          5349 => x"0c",
          5350 => x"76",
          5351 => x"38",
          5352 => x"11",
          5353 => x"81",
          5354 => x"51",
          5355 => x"13",
          5356 => x"8d",
          5357 => x"15",
          5358 => x"c5",
          5359 => x"90",
          5360 => x"0b",
          5361 => x"ff",
          5362 => x"15",
          5363 => x"2e",
          5364 => x"81",
          5365 => x"e4",
          5366 => x"88",
          5367 => x"ec",
          5368 => x"ff",
          5369 => x"81",
          5370 => x"06",
          5371 => x"81",
          5372 => x"51",
          5373 => x"82",
          5374 => x"80",
          5375 => x"85",
          5376 => x"15",
          5377 => x"14",
          5378 => x"3f",
          5379 => x"08",
          5380 => x"06",
          5381 => x"d4",
          5382 => x"81",
          5383 => x"38",
          5384 => x"d7",
          5385 => x"85",
          5386 => x"8b",
          5387 => x"2e",
          5388 => x"b3",
          5389 => x"14",
          5390 => x"3f",
          5391 => x"08",
          5392 => x"e4",
          5393 => x"81",
          5394 => x"84",
          5395 => x"d7",
          5396 => x"85",
          5397 => x"15",
          5398 => x"14",
          5399 => x"3f",
          5400 => x"08",
          5401 => x"76",
          5402 => x"9d",
          5403 => x"05",
          5404 => x"9d",
          5405 => x"86",
          5406 => x"0b",
          5407 => x"80",
          5408 => x"85",
          5409 => x"3d",
          5410 => x"3d",
          5411 => x"89",
          5412 => x"2e",
          5413 => x"08",
          5414 => x"2e",
          5415 => x"33",
          5416 => x"2e",
          5417 => x"13",
          5418 => x"22",
          5419 => x"76",
          5420 => x"06",
          5421 => x"13",
          5422 => x"92",
          5423 => x"ec",
          5424 => x"52",
          5425 => x"71",
          5426 => x"55",
          5427 => x"53",
          5428 => x"0c",
          5429 => x"85",
          5430 => x"3d",
          5431 => x"3d",
          5432 => x"05",
          5433 => x"89",
          5434 => x"52",
          5435 => x"3f",
          5436 => x"0b",
          5437 => x"08",
          5438 => x"82",
          5439 => x"82",
          5440 => x"90",
          5441 => x"55",
          5442 => x"2e",
          5443 => x"74",
          5444 => x"73",
          5445 => x"38",
          5446 => x"78",
          5447 => x"54",
          5448 => x"92",
          5449 => x"89",
          5450 => x"84",
          5451 => x"a9",
          5452 => x"ec",
          5453 => x"82",
          5454 => x"88",
          5455 => x"eb",
          5456 => x"02",
          5457 => x"e7",
          5458 => x"59",
          5459 => x"80",
          5460 => x"38",
          5461 => x"70",
          5462 => x"d0",
          5463 => x"3d",
          5464 => x"58",
          5465 => x"82",
          5466 => x"55",
          5467 => x"08",
          5468 => x"7a",
          5469 => x"8c",
          5470 => x"56",
          5471 => x"82",
          5472 => x"55",
          5473 => x"08",
          5474 => x"80",
          5475 => x"70",
          5476 => x"57",
          5477 => x"83",
          5478 => x"77",
          5479 => x"73",
          5480 => x"ab",
          5481 => x"2e",
          5482 => x"84",
          5483 => x"06",
          5484 => x"51",
          5485 => x"82",
          5486 => x"55",
          5487 => x"b2",
          5488 => x"06",
          5489 => x"b8",
          5490 => x"2a",
          5491 => x"51",
          5492 => x"2e",
          5493 => x"55",
          5494 => x"77",
          5495 => x"74",
          5496 => x"77",
          5497 => x"81",
          5498 => x"73",
          5499 => x"af",
          5500 => x"7a",
          5501 => x"3f",
          5502 => x"08",
          5503 => x"b2",
          5504 => x"8e",
          5505 => x"bc",
          5506 => x"a0",
          5507 => x"34",
          5508 => x"52",
          5509 => x"9e",
          5510 => x"62",
          5511 => x"d4",
          5512 => x"54",
          5513 => x"15",
          5514 => x"2e",
          5515 => x"7a",
          5516 => x"51",
          5517 => x"75",
          5518 => x"d4",
          5519 => x"97",
          5520 => x"ec",
          5521 => x"85",
          5522 => x"cc",
          5523 => x"74",
          5524 => x"02",
          5525 => x"70",
          5526 => x"81",
          5527 => x"56",
          5528 => x"86",
          5529 => x"82",
          5530 => x"81",
          5531 => x"06",
          5532 => x"80",
          5533 => x"75",
          5534 => x"73",
          5535 => x"38",
          5536 => x"94",
          5537 => x"7a",
          5538 => x"3f",
          5539 => x"08",
          5540 => x"8c",
          5541 => x"55",
          5542 => x"08",
          5543 => x"77",
          5544 => x"81",
          5545 => x"73",
          5546 => x"38",
          5547 => x"07",
          5548 => x"11",
          5549 => x"0c",
          5550 => x"0c",
          5551 => x"52",
          5552 => x"3f",
          5553 => x"08",
          5554 => x"08",
          5555 => x"63",
          5556 => x"5a",
          5557 => x"82",
          5558 => x"82",
          5559 => x"8c",
          5560 => x"7a",
          5561 => x"17",
          5562 => x"23",
          5563 => x"34",
          5564 => x"1a",
          5565 => x"9c",
          5566 => x"0b",
          5567 => x"77",
          5568 => x"81",
          5569 => x"73",
          5570 => x"8f",
          5571 => x"ec",
          5572 => x"81",
          5573 => x"85",
          5574 => x"1a",
          5575 => x"22",
          5576 => x"7b",
          5577 => x"a8",
          5578 => x"78",
          5579 => x"3f",
          5580 => x"08",
          5581 => x"ec",
          5582 => x"83",
          5583 => x"82",
          5584 => x"ff",
          5585 => x"06",
          5586 => x"55",
          5587 => x"56",
          5588 => x"05",
          5589 => x"80",
          5590 => x"77",
          5591 => x"38",
          5592 => x"06",
          5593 => x"c1",
          5594 => x"1a",
          5595 => x"38",
          5596 => x"06",
          5597 => x"2e",
          5598 => x"52",
          5599 => x"f6",
          5600 => x"ec",
          5601 => x"82",
          5602 => x"75",
          5603 => x"85",
          5604 => x"9c",
          5605 => x"39",
          5606 => x"74",
          5607 => x"85",
          5608 => x"3d",
          5609 => x"3d",
          5610 => x"65",
          5611 => x"5d",
          5612 => x"0c",
          5613 => x"05",
          5614 => x"f9",
          5615 => x"85",
          5616 => x"82",
          5617 => x"8a",
          5618 => x"33",
          5619 => x"2e",
          5620 => x"56",
          5621 => x"90",
          5622 => x"06",
          5623 => x"74",
          5624 => x"b6",
          5625 => x"82",
          5626 => x"34",
          5627 => x"aa",
          5628 => x"91",
          5629 => x"56",
          5630 => x"8c",
          5631 => x"1a",
          5632 => x"74",
          5633 => x"38",
          5634 => x"80",
          5635 => x"38",
          5636 => x"70",
          5637 => x"56",
          5638 => x"b2",
          5639 => x"11",
          5640 => x"77",
          5641 => x"5b",
          5642 => x"38",
          5643 => x"88",
          5644 => x"8f",
          5645 => x"08",
          5646 => x"d4",
          5647 => x"85",
          5648 => x"81",
          5649 => x"9f",
          5650 => x"2e",
          5651 => x"74",
          5652 => x"98",
          5653 => x"7e",
          5654 => x"3f",
          5655 => x"08",
          5656 => x"83",
          5657 => x"ec",
          5658 => x"89",
          5659 => x"77",
          5660 => x"d6",
          5661 => x"7f",
          5662 => x"58",
          5663 => x"75",
          5664 => x"75",
          5665 => x"77",
          5666 => x"7c",
          5667 => x"33",
          5668 => x"3f",
          5669 => x"08",
          5670 => x"7e",
          5671 => x"56",
          5672 => x"2e",
          5673 => x"16",
          5674 => x"55",
          5675 => x"94",
          5676 => x"53",
          5677 => x"b0",
          5678 => x"31",
          5679 => x"05",
          5680 => x"3f",
          5681 => x"56",
          5682 => x"9c",
          5683 => x"19",
          5684 => x"06",
          5685 => x"31",
          5686 => x"76",
          5687 => x"7b",
          5688 => x"08",
          5689 => x"d1",
          5690 => x"85",
          5691 => x"81",
          5692 => x"94",
          5693 => x"ff",
          5694 => x"05",
          5695 => x"ce",
          5696 => x"76",
          5697 => x"17",
          5698 => x"1e",
          5699 => x"18",
          5700 => x"5e",
          5701 => x"39",
          5702 => x"82",
          5703 => x"90",
          5704 => x"f2",
          5705 => x"63",
          5706 => x"40",
          5707 => x"7e",
          5708 => x"fc",
          5709 => x"51",
          5710 => x"82",
          5711 => x"55",
          5712 => x"08",
          5713 => x"18",
          5714 => x"80",
          5715 => x"74",
          5716 => x"39",
          5717 => x"70",
          5718 => x"81",
          5719 => x"56",
          5720 => x"80",
          5721 => x"38",
          5722 => x"0b",
          5723 => x"82",
          5724 => x"39",
          5725 => x"19",
          5726 => x"83",
          5727 => x"18",
          5728 => x"56",
          5729 => x"27",
          5730 => x"09",
          5731 => x"2e",
          5732 => x"94",
          5733 => x"83",
          5734 => x"56",
          5735 => x"38",
          5736 => x"22",
          5737 => x"89",
          5738 => x"55",
          5739 => x"75",
          5740 => x"18",
          5741 => x"9c",
          5742 => x"85",
          5743 => x"08",
          5744 => x"d7",
          5745 => x"85",
          5746 => x"82",
          5747 => x"80",
          5748 => x"38",
          5749 => x"ff",
          5750 => x"ff",
          5751 => x"38",
          5752 => x"0c",
          5753 => x"85",
          5754 => x"19",
          5755 => x"b0",
          5756 => x"19",
          5757 => x"81",
          5758 => x"74",
          5759 => x"3f",
          5760 => x"08",
          5761 => x"98",
          5762 => x"7e",
          5763 => x"3f",
          5764 => x"08",
          5765 => x"d2",
          5766 => x"ec",
          5767 => x"89",
          5768 => x"78",
          5769 => x"d5",
          5770 => x"7f",
          5771 => x"58",
          5772 => x"75",
          5773 => x"75",
          5774 => x"78",
          5775 => x"7c",
          5776 => x"33",
          5777 => x"3f",
          5778 => x"08",
          5779 => x"7e",
          5780 => x"78",
          5781 => x"74",
          5782 => x"38",
          5783 => x"b0",
          5784 => x"31",
          5785 => x"05",
          5786 => x"51",
          5787 => x"7e",
          5788 => x"83",
          5789 => x"89",
          5790 => x"db",
          5791 => x"08",
          5792 => x"26",
          5793 => x"51",
          5794 => x"82",
          5795 => x"fd",
          5796 => x"77",
          5797 => x"55",
          5798 => x"0c",
          5799 => x"83",
          5800 => x"80",
          5801 => x"55",
          5802 => x"83",
          5803 => x"9c",
          5804 => x"7e",
          5805 => x"3f",
          5806 => x"08",
          5807 => x"75",
          5808 => x"94",
          5809 => x"ff",
          5810 => x"05",
          5811 => x"3f",
          5812 => x"0b",
          5813 => x"7b",
          5814 => x"08",
          5815 => x"76",
          5816 => x"08",
          5817 => x"1c",
          5818 => x"08",
          5819 => x"5c",
          5820 => x"83",
          5821 => x"74",
          5822 => x"fd",
          5823 => x"18",
          5824 => x"07",
          5825 => x"19",
          5826 => x"75",
          5827 => x"0c",
          5828 => x"04",
          5829 => x"7a",
          5830 => x"05",
          5831 => x"56",
          5832 => x"82",
          5833 => x"57",
          5834 => x"08",
          5835 => x"90",
          5836 => x"86",
          5837 => x"06",
          5838 => x"73",
          5839 => x"e9",
          5840 => x"08",
          5841 => x"cc",
          5842 => x"85",
          5843 => x"82",
          5844 => x"80",
          5845 => x"16",
          5846 => x"33",
          5847 => x"55",
          5848 => x"34",
          5849 => x"53",
          5850 => x"08",
          5851 => x"3f",
          5852 => x"52",
          5853 => x"c9",
          5854 => x"88",
          5855 => x"96",
          5856 => x"c0",
          5857 => x"92",
          5858 => x"9a",
          5859 => x"81",
          5860 => x"34",
          5861 => x"af",
          5862 => x"ec",
          5863 => x"33",
          5864 => x"55",
          5865 => x"17",
          5866 => x"85",
          5867 => x"3d",
          5868 => x"3d",
          5869 => x"52",
          5870 => x"3f",
          5871 => x"08",
          5872 => x"ec",
          5873 => x"86",
          5874 => x"52",
          5875 => x"ba",
          5876 => x"ec",
          5877 => x"85",
          5878 => x"38",
          5879 => x"08",
          5880 => x"82",
          5881 => x"86",
          5882 => x"ff",
          5883 => x"3d",
          5884 => x"3f",
          5885 => x"0b",
          5886 => x"08",
          5887 => x"82",
          5888 => x"82",
          5889 => x"80",
          5890 => x"85",
          5891 => x"3d",
          5892 => x"3d",
          5893 => x"93",
          5894 => x"52",
          5895 => x"e9",
          5896 => x"85",
          5897 => x"82",
          5898 => x"80",
          5899 => x"58",
          5900 => x"3d",
          5901 => x"df",
          5902 => x"85",
          5903 => x"82",
          5904 => x"bc",
          5905 => x"c7",
          5906 => x"98",
          5907 => x"73",
          5908 => x"38",
          5909 => x"12",
          5910 => x"39",
          5911 => x"33",
          5912 => x"70",
          5913 => x"55",
          5914 => x"2e",
          5915 => x"7f",
          5916 => x"54",
          5917 => x"82",
          5918 => x"94",
          5919 => x"39",
          5920 => x"08",
          5921 => x"81",
          5922 => x"85",
          5923 => x"85",
          5924 => x"3d",
          5925 => x"3d",
          5926 => x"5b",
          5927 => x"34",
          5928 => x"3d",
          5929 => x"52",
          5930 => x"e8",
          5931 => x"85",
          5932 => x"82",
          5933 => x"82",
          5934 => x"43",
          5935 => x"11",
          5936 => x"58",
          5937 => x"80",
          5938 => x"38",
          5939 => x"3d",
          5940 => x"d5",
          5941 => x"85",
          5942 => x"82",
          5943 => x"82",
          5944 => x"52",
          5945 => x"98",
          5946 => x"ec",
          5947 => x"85",
          5948 => x"c0",
          5949 => x"7b",
          5950 => x"3f",
          5951 => x"08",
          5952 => x"74",
          5953 => x"3f",
          5954 => x"08",
          5955 => x"ec",
          5956 => x"38",
          5957 => x"51",
          5958 => x"82",
          5959 => x"57",
          5960 => x"08",
          5961 => x"52",
          5962 => x"d1",
          5963 => x"85",
          5964 => x"a6",
          5965 => x"74",
          5966 => x"3f",
          5967 => x"08",
          5968 => x"ec",
          5969 => x"cc",
          5970 => x"2e",
          5971 => x"86",
          5972 => x"81",
          5973 => x"81",
          5974 => x"3d",
          5975 => x"52",
          5976 => x"a8",
          5977 => x"3d",
          5978 => x"11",
          5979 => x"5a",
          5980 => x"2e",
          5981 => x"b9",
          5982 => x"16",
          5983 => x"33",
          5984 => x"73",
          5985 => x"16",
          5986 => x"26",
          5987 => x"75",
          5988 => x"38",
          5989 => x"05",
          5990 => x"6f",
          5991 => x"ff",
          5992 => x"55",
          5993 => x"74",
          5994 => x"38",
          5995 => x"11",
          5996 => x"74",
          5997 => x"39",
          5998 => x"09",
          5999 => x"38",
          6000 => x"11",
          6001 => x"74",
          6002 => x"82",
          6003 => x"70",
          6004 => x"ff",
          6005 => x"70",
          6006 => x"56",
          6007 => x"76",
          6008 => x"81",
          6009 => x"70",
          6010 => x"56",
          6011 => x"82",
          6012 => x"78",
          6013 => x"80",
          6014 => x"27",
          6015 => x"19",
          6016 => x"7a",
          6017 => x"5c",
          6018 => x"55",
          6019 => x"7a",
          6020 => x"5c",
          6021 => x"2e",
          6022 => x"85",
          6023 => x"94",
          6024 => x"81",
          6025 => x"73",
          6026 => x"81",
          6027 => x"7a",
          6028 => x"38",
          6029 => x"76",
          6030 => x"0c",
          6031 => x"04",
          6032 => x"7b",
          6033 => x"fc",
          6034 => x"53",
          6035 => x"ba",
          6036 => x"ec",
          6037 => x"85",
          6038 => x"fc",
          6039 => x"33",
          6040 => x"f4",
          6041 => x"08",
          6042 => x"27",
          6043 => x"15",
          6044 => x"2a",
          6045 => x"51",
          6046 => x"83",
          6047 => x"94",
          6048 => x"80",
          6049 => x"0c",
          6050 => x"2e",
          6051 => x"79",
          6052 => x"70",
          6053 => x"51",
          6054 => x"2e",
          6055 => x"52",
          6056 => x"fe",
          6057 => x"82",
          6058 => x"ff",
          6059 => x"70",
          6060 => x"fe",
          6061 => x"82",
          6062 => x"73",
          6063 => x"76",
          6064 => x"70",
          6065 => x"94",
          6066 => x"71",
          6067 => x"08",
          6068 => x"53",
          6069 => x"15",
          6070 => x"a6",
          6071 => x"74",
          6072 => x"3f",
          6073 => x"08",
          6074 => x"ec",
          6075 => x"81",
          6076 => x"85",
          6077 => x"2e",
          6078 => x"82",
          6079 => x"88",
          6080 => x"98",
          6081 => x"80",
          6082 => x"38",
          6083 => x"80",
          6084 => x"77",
          6085 => x"08",
          6086 => x"0c",
          6087 => x"70",
          6088 => x"81",
          6089 => x"5a",
          6090 => x"2e",
          6091 => x"52",
          6092 => x"cf",
          6093 => x"ec",
          6094 => x"85",
          6095 => x"38",
          6096 => x"08",
          6097 => x"73",
          6098 => x"c6",
          6099 => x"85",
          6100 => x"73",
          6101 => x"38",
          6102 => x"af",
          6103 => x"73",
          6104 => x"27",
          6105 => x"98",
          6106 => x"a0",
          6107 => x"08",
          6108 => x"0c",
          6109 => x"06",
          6110 => x"2e",
          6111 => x"52",
          6112 => x"f2",
          6113 => x"ec",
          6114 => x"82",
          6115 => x"34",
          6116 => x"c4",
          6117 => x"91",
          6118 => x"53",
          6119 => x"89",
          6120 => x"ec",
          6121 => x"94",
          6122 => x"8c",
          6123 => x"27",
          6124 => x"8c",
          6125 => x"15",
          6126 => x"07",
          6127 => x"16",
          6128 => x"ff",
          6129 => x"80",
          6130 => x"77",
          6131 => x"2e",
          6132 => x"9c",
          6133 => x"53",
          6134 => x"ec",
          6135 => x"0d",
          6136 => x"0d",
          6137 => x"54",
          6138 => x"81",
          6139 => x"53",
          6140 => x"05",
          6141 => x"84",
          6142 => x"dd",
          6143 => x"ec",
          6144 => x"85",
          6145 => x"ea",
          6146 => x"0c",
          6147 => x"51",
          6148 => x"82",
          6149 => x"55",
          6150 => x"08",
          6151 => x"ab",
          6152 => x"98",
          6153 => x"80",
          6154 => x"38",
          6155 => x"70",
          6156 => x"81",
          6157 => x"57",
          6158 => x"ad",
          6159 => x"08",
          6160 => x"d3",
          6161 => x"85",
          6162 => x"17",
          6163 => x"86",
          6164 => x"17",
          6165 => x"75",
          6166 => x"3f",
          6167 => x"08",
          6168 => x"2e",
          6169 => x"85",
          6170 => x"86",
          6171 => x"2e",
          6172 => x"76",
          6173 => x"73",
          6174 => x"0c",
          6175 => x"04",
          6176 => x"76",
          6177 => x"05",
          6178 => x"53",
          6179 => x"82",
          6180 => x"87",
          6181 => x"ec",
          6182 => x"86",
          6183 => x"fb",
          6184 => x"79",
          6185 => x"05",
          6186 => x"56",
          6187 => x"3f",
          6188 => x"08",
          6189 => x"ec",
          6190 => x"38",
          6191 => x"82",
          6192 => x"52",
          6193 => x"d6",
          6194 => x"ec",
          6195 => x"cc",
          6196 => x"ec",
          6197 => x"51",
          6198 => x"82",
          6199 => x"53",
          6200 => x"08",
          6201 => x"81",
          6202 => x"80",
          6203 => x"82",
          6204 => x"a8",
          6205 => x"73",
          6206 => x"3f",
          6207 => x"51",
          6208 => x"82",
          6209 => x"84",
          6210 => x"81",
          6211 => x"07",
          6212 => x"82",
          6213 => x"06",
          6214 => x"54",
          6215 => x"ec",
          6216 => x"0d",
          6217 => x"0d",
          6218 => x"53",
          6219 => x"53",
          6220 => x"56",
          6221 => x"82",
          6222 => x"55",
          6223 => x"08",
          6224 => x"52",
          6225 => x"dd",
          6226 => x"ec",
          6227 => x"85",
          6228 => x"38",
          6229 => x"05",
          6230 => x"2b",
          6231 => x"80",
          6232 => x"86",
          6233 => x"76",
          6234 => x"38",
          6235 => x"51",
          6236 => x"74",
          6237 => x"0c",
          6238 => x"04",
          6239 => x"63",
          6240 => x"80",
          6241 => x"ec",
          6242 => x"3d",
          6243 => x"3f",
          6244 => x"08",
          6245 => x"ec",
          6246 => x"38",
          6247 => x"73",
          6248 => x"08",
          6249 => x"13",
          6250 => x"58",
          6251 => x"26",
          6252 => x"7c",
          6253 => x"39",
          6254 => x"d3",
          6255 => x"81",
          6256 => x"85",
          6257 => x"33",
          6258 => x"81",
          6259 => x"06",
          6260 => x"82",
          6261 => x"76",
          6262 => x"f0",
          6263 => x"c7",
          6264 => x"ec",
          6265 => x"d0",
          6266 => x"ec",
          6267 => x"cd",
          6268 => x"ec",
          6269 => x"05",
          6270 => x"ec",
          6271 => x"25",
          6272 => x"19",
          6273 => x"5a",
          6274 => x"08",
          6275 => x"38",
          6276 => x"a4",
          6277 => x"85",
          6278 => x"58",
          6279 => x"77",
          6280 => x"7d",
          6281 => x"be",
          6282 => x"85",
          6283 => x"82",
          6284 => x"80",
          6285 => x"70",
          6286 => x"ff",
          6287 => x"56",
          6288 => x"2e",
          6289 => x"a0",
          6290 => x"51",
          6291 => x"3f",
          6292 => x"08",
          6293 => x"06",
          6294 => x"05",
          6295 => x"1b",
          6296 => x"5b",
          6297 => x"39",
          6298 => x"ff",
          6299 => x"82",
          6300 => x"f0",
          6301 => x"09",
          6302 => x"80",
          6303 => x"19",
          6304 => x"54",
          6305 => x"06",
          6306 => x"79",
          6307 => x"78",
          6308 => x"79",
          6309 => x"84",
          6310 => x"07",
          6311 => x"84",
          6312 => x"82",
          6313 => x"92",
          6314 => x"f9",
          6315 => x"8a",
          6316 => x"53",
          6317 => x"e3",
          6318 => x"85",
          6319 => x"82",
          6320 => x"81",
          6321 => x"17",
          6322 => x"81",
          6323 => x"17",
          6324 => x"2a",
          6325 => x"51",
          6326 => x"55",
          6327 => x"81",
          6328 => x"17",
          6329 => x"8c",
          6330 => x"81",
          6331 => x"9b",
          6332 => x"ec",
          6333 => x"17",
          6334 => x"51",
          6335 => x"82",
          6336 => x"74",
          6337 => x"56",
          6338 => x"98",
          6339 => x"76",
          6340 => x"93",
          6341 => x"ec",
          6342 => x"09",
          6343 => x"38",
          6344 => x"85",
          6345 => x"2e",
          6346 => x"85",
          6347 => x"a3",
          6348 => x"38",
          6349 => x"85",
          6350 => x"15",
          6351 => x"38",
          6352 => x"53",
          6353 => x"08",
          6354 => x"c3",
          6355 => x"85",
          6356 => x"94",
          6357 => x"18",
          6358 => x"33",
          6359 => x"54",
          6360 => x"34",
          6361 => x"85",
          6362 => x"18",
          6363 => x"74",
          6364 => x"0c",
          6365 => x"04",
          6366 => x"82",
          6367 => x"ff",
          6368 => x"a1",
          6369 => x"d1",
          6370 => x"ec",
          6371 => x"85",
          6372 => x"f7",
          6373 => x"a1",
          6374 => x"95",
          6375 => x"58",
          6376 => x"82",
          6377 => x"55",
          6378 => x"08",
          6379 => x"02",
          6380 => x"33",
          6381 => x"70",
          6382 => x"55",
          6383 => x"73",
          6384 => x"75",
          6385 => x"80",
          6386 => x"bf",
          6387 => x"d6",
          6388 => x"81",
          6389 => x"87",
          6390 => x"af",
          6391 => x"78",
          6392 => x"3f",
          6393 => x"08",
          6394 => x"70",
          6395 => x"55",
          6396 => x"2e",
          6397 => x"78",
          6398 => x"ec",
          6399 => x"08",
          6400 => x"38",
          6401 => x"85",
          6402 => x"76",
          6403 => x"70",
          6404 => x"8a",
          6405 => x"ec",
          6406 => x"85",
          6407 => x"eb",
          6408 => x"ec",
          6409 => x"51",
          6410 => x"82",
          6411 => x"55",
          6412 => x"08",
          6413 => x"55",
          6414 => x"82",
          6415 => x"84",
          6416 => x"82",
          6417 => x"80",
          6418 => x"51",
          6419 => x"82",
          6420 => x"82",
          6421 => x"09",
          6422 => x"82",
          6423 => x"07",
          6424 => x"55",
          6425 => x"2e",
          6426 => x"80",
          6427 => x"80",
          6428 => x"77",
          6429 => x"3f",
          6430 => x"08",
          6431 => x"38",
          6432 => x"ba",
          6433 => x"85",
          6434 => x"74",
          6435 => x"0c",
          6436 => x"04",
          6437 => x"82",
          6438 => x"c0",
          6439 => x"3d",
          6440 => x"3f",
          6441 => x"08",
          6442 => x"ec",
          6443 => x"38",
          6444 => x"52",
          6445 => x"52",
          6446 => x"3f",
          6447 => x"08",
          6448 => x"ec",
          6449 => x"88",
          6450 => x"39",
          6451 => x"08",
          6452 => x"81",
          6453 => x"38",
          6454 => x"05",
          6455 => x"2a",
          6456 => x"55",
          6457 => x"81",
          6458 => x"5a",
          6459 => x"3d",
          6460 => x"c1",
          6461 => x"85",
          6462 => x"55",
          6463 => x"ec",
          6464 => x"87",
          6465 => x"ec",
          6466 => x"09",
          6467 => x"38",
          6468 => x"85",
          6469 => x"2e",
          6470 => x"86",
          6471 => x"81",
          6472 => x"81",
          6473 => x"85",
          6474 => x"78",
          6475 => x"3f",
          6476 => x"08",
          6477 => x"ec",
          6478 => x"38",
          6479 => x"52",
          6480 => x"ff",
          6481 => x"78",
          6482 => x"b4",
          6483 => x"54",
          6484 => x"15",
          6485 => x"b2",
          6486 => x"ca",
          6487 => x"b5",
          6488 => x"53",
          6489 => x"53",
          6490 => x"3f",
          6491 => x"b4",
          6492 => x"d4",
          6493 => x"b5",
          6494 => x"54",
          6495 => x"d5",
          6496 => x"53",
          6497 => x"11",
          6498 => x"aa",
          6499 => x"81",
          6500 => x"34",
          6501 => x"f7",
          6502 => x"ec",
          6503 => x"85",
          6504 => x"38",
          6505 => x"0a",
          6506 => x"05",
          6507 => x"94",
          6508 => x"64",
          6509 => x"c8",
          6510 => x"54",
          6511 => x"15",
          6512 => x"81",
          6513 => x"34",
          6514 => x"b7",
          6515 => x"85",
          6516 => x"8b",
          6517 => x"75",
          6518 => x"ff",
          6519 => x"73",
          6520 => x"0c",
          6521 => x"04",
          6522 => x"a9",
          6523 => x"51",
          6524 => x"82",
          6525 => x"ff",
          6526 => x"a9",
          6527 => x"d9",
          6528 => x"ec",
          6529 => x"85",
          6530 => x"d3",
          6531 => x"a9",
          6532 => x"9d",
          6533 => x"58",
          6534 => x"82",
          6535 => x"55",
          6536 => x"08",
          6537 => x"02",
          6538 => x"33",
          6539 => x"54",
          6540 => x"82",
          6541 => x"53",
          6542 => x"52",
          6543 => x"88",
          6544 => x"b4",
          6545 => x"53",
          6546 => x"3d",
          6547 => x"ff",
          6548 => x"aa",
          6549 => x"73",
          6550 => x"3f",
          6551 => x"08",
          6552 => x"ec",
          6553 => x"63",
          6554 => x"81",
          6555 => x"65",
          6556 => x"2e",
          6557 => x"55",
          6558 => x"82",
          6559 => x"84",
          6560 => x"06",
          6561 => x"73",
          6562 => x"3f",
          6563 => x"08",
          6564 => x"ec",
          6565 => x"38",
          6566 => x"53",
          6567 => x"95",
          6568 => x"16",
          6569 => x"cb",
          6570 => x"05",
          6571 => x"34",
          6572 => x"70",
          6573 => x"81",
          6574 => x"55",
          6575 => x"74",
          6576 => x"73",
          6577 => x"78",
          6578 => x"83",
          6579 => x"16",
          6580 => x"2a",
          6581 => x"51",
          6582 => x"80",
          6583 => x"38",
          6584 => x"80",
          6585 => x"52",
          6586 => x"91",
          6587 => x"ec",
          6588 => x"51",
          6589 => x"3f",
          6590 => x"85",
          6591 => x"2e",
          6592 => x"82",
          6593 => x"52",
          6594 => x"b4",
          6595 => x"85",
          6596 => x"80",
          6597 => x"58",
          6598 => x"ec",
          6599 => x"38",
          6600 => x"54",
          6601 => x"09",
          6602 => x"38",
          6603 => x"52",
          6604 => x"82",
          6605 => x"81",
          6606 => x"34",
          6607 => x"85",
          6608 => x"38",
          6609 => x"9d",
          6610 => x"ec",
          6611 => x"85",
          6612 => x"38",
          6613 => x"b4",
          6614 => x"85",
          6615 => x"74",
          6616 => x"0c",
          6617 => x"04",
          6618 => x"02",
          6619 => x"33",
          6620 => x"80",
          6621 => x"57",
          6622 => x"95",
          6623 => x"52",
          6624 => x"d2",
          6625 => x"85",
          6626 => x"82",
          6627 => x"80",
          6628 => x"5a",
          6629 => x"3d",
          6630 => x"c9",
          6631 => x"85",
          6632 => x"82",
          6633 => x"b8",
          6634 => x"cf",
          6635 => x"a0",
          6636 => x"55",
          6637 => x"75",
          6638 => x"71",
          6639 => x"33",
          6640 => x"74",
          6641 => x"57",
          6642 => x"8b",
          6643 => x"54",
          6644 => x"15",
          6645 => x"ff",
          6646 => x"82",
          6647 => x"55",
          6648 => x"ec",
          6649 => x"0d",
          6650 => x"0d",
          6651 => x"53",
          6652 => x"05",
          6653 => x"51",
          6654 => x"82",
          6655 => x"55",
          6656 => x"08",
          6657 => x"76",
          6658 => x"93",
          6659 => x"51",
          6660 => x"82",
          6661 => x"55",
          6662 => x"08",
          6663 => x"80",
          6664 => x"81",
          6665 => x"86",
          6666 => x"38",
          6667 => x"86",
          6668 => x"90",
          6669 => x"54",
          6670 => x"ff",
          6671 => x"76",
          6672 => x"83",
          6673 => x"51",
          6674 => x"3f",
          6675 => x"08",
          6676 => x"85",
          6677 => x"3d",
          6678 => x"3d",
          6679 => x"5c",
          6680 => x"98",
          6681 => x"52",
          6682 => x"d0",
          6683 => x"85",
          6684 => x"85",
          6685 => x"81",
          6686 => x"85",
          6687 => x"80",
          6688 => x"57",
          6689 => x"81",
          6690 => x"70",
          6691 => x"55",
          6692 => x"80",
          6693 => x"5d",
          6694 => x"52",
          6695 => x"52",
          6696 => x"fa",
          6697 => x"ec",
          6698 => x"85",
          6699 => x"d1",
          6700 => x"73",
          6701 => x"3f",
          6702 => x"08",
          6703 => x"ec",
          6704 => x"82",
          6705 => x"82",
          6706 => x"65",
          6707 => x"78",
          6708 => x"7b",
          6709 => x"55",
          6710 => x"34",
          6711 => x"8a",
          6712 => x"38",
          6713 => x"1a",
          6714 => x"34",
          6715 => x"9e",
          6716 => x"70",
          6717 => x"51",
          6718 => x"a0",
          6719 => x"8e",
          6720 => x"2e",
          6721 => x"86",
          6722 => x"34",
          6723 => x"09",
          6724 => x"78",
          6725 => x"51",
          6726 => x"2e",
          6727 => x"73",
          6728 => x"38",
          6729 => x"08",
          6730 => x"b0",
          6731 => x"85",
          6732 => x"82",
          6733 => x"a7",
          6734 => x"33",
          6735 => x"c3",
          6736 => x"2e",
          6737 => x"e4",
          6738 => x"2e",
          6739 => x"56",
          6740 => x"05",
          6741 => x"a3",
          6742 => x"ec",
          6743 => x"76",
          6744 => x"0c",
          6745 => x"04",
          6746 => x"82",
          6747 => x"ff",
          6748 => x"9d",
          6749 => x"e1",
          6750 => x"ec",
          6751 => x"ec",
          6752 => x"82",
          6753 => x"83",
          6754 => x"53",
          6755 => x"3d",
          6756 => x"ff",
          6757 => x"73",
          6758 => x"70",
          6759 => x"52",
          6760 => x"9f",
          6761 => x"bc",
          6762 => x"74",
          6763 => x"6d",
          6764 => x"70",
          6765 => x"ae",
          6766 => x"85",
          6767 => x"2e",
          6768 => x"70",
          6769 => x"57",
          6770 => x"bd",
          6771 => x"ec",
          6772 => x"8d",
          6773 => x"2b",
          6774 => x"81",
          6775 => x"86",
          6776 => x"ec",
          6777 => x"9f",
          6778 => x"ff",
          6779 => x"54",
          6780 => x"8a",
          6781 => x"70",
          6782 => x"06",
          6783 => x"ff",
          6784 => x"38",
          6785 => x"15",
          6786 => x"80",
          6787 => x"74",
          6788 => x"b4",
          6789 => x"c9",
          6790 => x"ec",
          6791 => x"81",
          6792 => x"88",
          6793 => x"26",
          6794 => x"39",
          6795 => x"86",
          6796 => x"81",
          6797 => x"ff",
          6798 => x"38",
          6799 => x"54",
          6800 => x"81",
          6801 => x"81",
          6802 => x"78",
          6803 => x"5a",
          6804 => x"6d",
          6805 => x"81",
          6806 => x"57",
          6807 => x"9f",
          6808 => x"38",
          6809 => x"54",
          6810 => x"81",
          6811 => x"b1",
          6812 => x"2e",
          6813 => x"a7",
          6814 => x"15",
          6815 => x"54",
          6816 => x"09",
          6817 => x"38",
          6818 => x"76",
          6819 => x"41",
          6820 => x"52",
          6821 => x"52",
          6822 => x"82",
          6823 => x"ec",
          6824 => x"85",
          6825 => x"f7",
          6826 => x"74",
          6827 => x"b4",
          6828 => x"ec",
          6829 => x"85",
          6830 => x"38",
          6831 => x"38",
          6832 => x"74",
          6833 => x"39",
          6834 => x"08",
          6835 => x"81",
          6836 => x"38",
          6837 => x"74",
          6838 => x"38",
          6839 => x"51",
          6840 => x"3f",
          6841 => x"08",
          6842 => x"ec",
          6843 => x"a0",
          6844 => x"ec",
          6845 => x"51",
          6846 => x"3f",
          6847 => x"0b",
          6848 => x"8b",
          6849 => x"67",
          6850 => x"e7",
          6851 => x"81",
          6852 => x"34",
          6853 => x"ad",
          6854 => x"85",
          6855 => x"73",
          6856 => x"85",
          6857 => x"3d",
          6858 => x"3d",
          6859 => x"02",
          6860 => x"cb",
          6861 => x"3d",
          6862 => x"72",
          6863 => x"5a",
          6864 => x"82",
          6865 => x"58",
          6866 => x"08",
          6867 => x"91",
          6868 => x"77",
          6869 => x"7c",
          6870 => x"38",
          6871 => x"59",
          6872 => x"90",
          6873 => x"81",
          6874 => x"06",
          6875 => x"73",
          6876 => x"54",
          6877 => x"82",
          6878 => x"39",
          6879 => x"8d",
          6880 => x"11",
          6881 => x"2b",
          6882 => x"54",
          6883 => x"fe",
          6884 => x"ff",
          6885 => x"70",
          6886 => x"70",
          6887 => x"2a",
          6888 => x"08",
          6889 => x"08",
          6890 => x"5d",
          6891 => x"77",
          6892 => x"98",
          6893 => x"26",
          6894 => x"57",
          6895 => x"59",
          6896 => x"52",
          6897 => x"ad",
          6898 => x"15",
          6899 => x"98",
          6900 => x"26",
          6901 => x"55",
          6902 => x"08",
          6903 => x"97",
          6904 => x"ec",
          6905 => x"ff",
          6906 => x"85",
          6907 => x"38",
          6908 => x"75",
          6909 => x"81",
          6910 => x"93",
          6911 => x"80",
          6912 => x"2e",
          6913 => x"ff",
          6914 => x"58",
          6915 => x"7d",
          6916 => x"38",
          6917 => x"55",
          6918 => x"b4",
          6919 => x"56",
          6920 => x"09",
          6921 => x"38",
          6922 => x"53",
          6923 => x"51",
          6924 => x"3f",
          6925 => x"08",
          6926 => x"ec",
          6927 => x"38",
          6928 => x"ff",
          6929 => x"5c",
          6930 => x"84",
          6931 => x"5c",
          6932 => x"12",
          6933 => x"80",
          6934 => x"78",
          6935 => x"7c",
          6936 => x"90",
          6937 => x"c0",
          6938 => x"90",
          6939 => x"15",
          6940 => x"90",
          6941 => x"54",
          6942 => x"91",
          6943 => x"31",
          6944 => x"84",
          6945 => x"07",
          6946 => x"16",
          6947 => x"73",
          6948 => x"0c",
          6949 => x"04",
          6950 => x"6b",
          6951 => x"05",
          6952 => x"33",
          6953 => x"5a",
          6954 => x"9a",
          6955 => x"80",
          6956 => x"ec",
          6957 => x"82",
          6958 => x"ec",
          6959 => x"82",
          6960 => x"08",
          6961 => x"80",
          6962 => x"80",
          6963 => x"85",
          6964 => x"ff",
          6965 => x"52",
          6966 => x"a0",
          6967 => x"85",
          6968 => x"ff",
          6969 => x"06",
          6970 => x"56",
          6971 => x"38",
          6972 => x"70",
          6973 => x"55",
          6974 => x"8b",
          6975 => x"3d",
          6976 => x"83",
          6977 => x"ff",
          6978 => x"82",
          6979 => x"99",
          6980 => x"74",
          6981 => x"38",
          6982 => x"80",
          6983 => x"ff",
          6984 => x"55",
          6985 => x"83",
          6986 => x"78",
          6987 => x"38",
          6988 => x"26",
          6989 => x"81",
          6990 => x"8b",
          6991 => x"79",
          6992 => x"80",
          6993 => x"93",
          6994 => x"39",
          6995 => x"6e",
          6996 => x"89",
          6997 => x"48",
          6998 => x"83",
          6999 => x"61",
          7000 => x"70",
          7001 => x"07",
          7002 => x"56",
          7003 => x"38",
          7004 => x"05",
          7005 => x"7e",
          7006 => x"bd",
          7007 => x"82",
          7008 => x"8a",
          7009 => x"83",
          7010 => x"06",
          7011 => x"08",
          7012 => x"74",
          7013 => x"41",
          7014 => x"56",
          7015 => x"8a",
          7016 => x"61",
          7017 => x"55",
          7018 => x"27",
          7019 => x"93",
          7020 => x"80",
          7021 => x"38",
          7022 => x"70",
          7023 => x"43",
          7024 => x"95",
          7025 => x"06",
          7026 => x"2e",
          7027 => x"77",
          7028 => x"74",
          7029 => x"8a",
          7030 => x"06",
          7031 => x"82",
          7032 => x"2e",
          7033 => x"78",
          7034 => x"2e",
          7035 => x"80",
          7036 => x"ae",
          7037 => x"2a",
          7038 => x"82",
          7039 => x"56",
          7040 => x"2e",
          7041 => x"77",
          7042 => x"82",
          7043 => x"79",
          7044 => x"70",
          7045 => x"5a",
          7046 => x"86",
          7047 => x"27",
          7048 => x"52",
          7049 => x"c1",
          7050 => x"85",
          7051 => x"2b",
          7052 => x"89",
          7053 => x"a0",
          7054 => x"82",
          7055 => x"fc",
          7056 => x"56",
          7057 => x"f0",
          7058 => x"80",
          7059 => x"dd",
          7060 => x"38",
          7061 => x"57",
          7062 => x"80",
          7063 => x"5a",
          7064 => x"9d",
          7065 => x"26",
          7066 => x"80",
          7067 => x"10",
          7068 => x"22",
          7069 => x"74",
          7070 => x"38",
          7071 => x"ee",
          7072 => x"66",
          7073 => x"85",
          7074 => x"ec",
          7075 => x"ec",
          7076 => x"05",
          7077 => x"ec",
          7078 => x"26",
          7079 => x"0b",
          7080 => x"08",
          7081 => x"85",
          7082 => x"12",
          7083 => x"83",
          7084 => x"56",
          7085 => x"17",
          7086 => x"81",
          7087 => x"60",
          7088 => x"65",
          7089 => x"12",
          7090 => x"09",
          7091 => x"72",
          7092 => x"5c",
          7093 => x"59",
          7094 => x"2e",
          7095 => x"89",
          7096 => x"60",
          7097 => x"84",
          7098 => x"5d",
          7099 => x"70",
          7100 => x"68",
          7101 => x"74",
          7102 => x"b1",
          7103 => x"31",
          7104 => x"53",
          7105 => x"52",
          7106 => x"81",
          7107 => x"ec",
          7108 => x"83",
          7109 => x"06",
          7110 => x"85",
          7111 => x"ff",
          7112 => x"dd",
          7113 => x"85",
          7114 => x"2a",
          7115 => x"b7",
          7116 => x"39",
          7117 => x"09",
          7118 => x"c5",
          7119 => x"f5",
          7120 => x"ec",
          7121 => x"38",
          7122 => x"79",
          7123 => x"80",
          7124 => x"38",
          7125 => x"8f",
          7126 => x"06",
          7127 => x"2e",
          7128 => x"5e",
          7129 => x"82",
          7130 => x"9f",
          7131 => x"38",
          7132 => x"38",
          7133 => x"81",
          7134 => x"fc",
          7135 => x"ad",
          7136 => x"7d",
          7137 => x"81",
          7138 => x"7d",
          7139 => x"78",
          7140 => x"74",
          7141 => x"8e",
          7142 => x"9e",
          7143 => x"53",
          7144 => x"51",
          7145 => x"3f",
          7146 => x"fe",
          7147 => x"51",
          7148 => x"3f",
          7149 => x"8b",
          7150 => x"a0",
          7151 => x"8d",
          7152 => x"83",
          7153 => x"52",
          7154 => x"ff",
          7155 => x"81",
          7156 => x"34",
          7157 => x"70",
          7158 => x"70",
          7159 => x"80",
          7160 => x"55",
          7161 => x"ff",
          7162 => x"66",
          7163 => x"ff",
          7164 => x"38",
          7165 => x"ff",
          7166 => x"1b",
          7167 => x"a6",
          7168 => x"74",
          7169 => x"51",
          7170 => x"3f",
          7171 => x"1c",
          7172 => x"98",
          7173 => x"a0",
          7174 => x"ff",
          7175 => x"51",
          7176 => x"3f",
          7177 => x"1b",
          7178 => x"98",
          7179 => x"2e",
          7180 => x"80",
          7181 => x"88",
          7182 => x"80",
          7183 => x"ff",
          7184 => x"7c",
          7185 => x"51",
          7186 => x"3f",
          7187 => x"1b",
          7188 => x"f0",
          7189 => x"b0",
          7190 => x"9f",
          7191 => x"52",
          7192 => x"ff",
          7193 => x"ff",
          7194 => x"c0",
          7195 => x"0b",
          7196 => x"34",
          7197 => x"fe",
          7198 => x"c7",
          7199 => x"39",
          7200 => x"0a",
          7201 => x"51",
          7202 => x"3f",
          7203 => x"ff",
          7204 => x"1b",
          7205 => x"8e",
          7206 => x"0b",
          7207 => x"a9",
          7208 => x"34",
          7209 => x"ff",
          7210 => x"1b",
          7211 => x"c3",
          7212 => x"d5",
          7213 => x"1b",
          7214 => x"ff",
          7215 => x"81",
          7216 => x"7a",
          7217 => x"ff",
          7218 => x"81",
          7219 => x"ec",
          7220 => x"38",
          7221 => x"09",
          7222 => x"ee",
          7223 => x"60",
          7224 => x"7a",
          7225 => x"ff",
          7226 => x"84",
          7227 => x"52",
          7228 => x"9f",
          7229 => x"8b",
          7230 => x"52",
          7231 => x"9e",
          7232 => x"8a",
          7233 => x"52",
          7234 => x"51",
          7235 => x"3f",
          7236 => x"83",
          7237 => x"ff",
          7238 => x"82",
          7239 => x"1b",
          7240 => x"a0",
          7241 => x"d5",
          7242 => x"ff",
          7243 => x"75",
          7244 => x"05",
          7245 => x"7e",
          7246 => x"99",
          7247 => x"60",
          7248 => x"52",
          7249 => x"9a",
          7250 => x"53",
          7251 => x"51",
          7252 => x"3f",
          7253 => x"58",
          7254 => x"09",
          7255 => x"38",
          7256 => x"51",
          7257 => x"3f",
          7258 => x"1b",
          7259 => x"d4",
          7260 => x"52",
          7261 => x"91",
          7262 => x"ff",
          7263 => x"81",
          7264 => x"f8",
          7265 => x"7a",
          7266 => x"b8",
          7267 => x"61",
          7268 => x"26",
          7269 => x"57",
          7270 => x"53",
          7271 => x"51",
          7272 => x"3f",
          7273 => x"08",
          7274 => x"84",
          7275 => x"85",
          7276 => x"7a",
          7277 => x"de",
          7278 => x"75",
          7279 => x"56",
          7280 => x"81",
          7281 => x"80",
          7282 => x"38",
          7283 => x"83",
          7284 => x"63",
          7285 => x"74",
          7286 => x"38",
          7287 => x"54",
          7288 => x"52",
          7289 => x"98",
          7290 => x"85",
          7291 => x"c1",
          7292 => x"75",
          7293 => x"56",
          7294 => x"8c",
          7295 => x"2e",
          7296 => x"56",
          7297 => x"ff",
          7298 => x"84",
          7299 => x"2e",
          7300 => x"56",
          7301 => x"58",
          7302 => x"38",
          7303 => x"77",
          7304 => x"ff",
          7305 => x"82",
          7306 => x"78",
          7307 => x"f6",
          7308 => x"1b",
          7309 => x"34",
          7310 => x"16",
          7311 => x"82",
          7312 => x"83",
          7313 => x"84",
          7314 => x"67",
          7315 => x"fd",
          7316 => x"51",
          7317 => x"3f",
          7318 => x"16",
          7319 => x"ec",
          7320 => x"bf",
          7321 => x"86",
          7322 => x"85",
          7323 => x"16",
          7324 => x"83",
          7325 => x"ff",
          7326 => x"66",
          7327 => x"1b",
          7328 => x"c0",
          7329 => x"77",
          7330 => x"7e",
          7331 => x"c5",
          7332 => x"82",
          7333 => x"a2",
          7334 => x"80",
          7335 => x"ff",
          7336 => x"81",
          7337 => x"ec",
          7338 => x"89",
          7339 => x"8a",
          7340 => x"86",
          7341 => x"ec",
          7342 => x"82",
          7343 => x"99",
          7344 => x"f5",
          7345 => x"60",
          7346 => x"79",
          7347 => x"5a",
          7348 => x"78",
          7349 => x"8d",
          7350 => x"55",
          7351 => x"fc",
          7352 => x"51",
          7353 => x"7a",
          7354 => x"81",
          7355 => x"8c",
          7356 => x"74",
          7357 => x"38",
          7358 => x"81",
          7359 => x"81",
          7360 => x"8a",
          7361 => x"06",
          7362 => x"76",
          7363 => x"76",
          7364 => x"55",
          7365 => x"ec",
          7366 => x"0d",
          7367 => x"0d",
          7368 => x"05",
          7369 => x"59",
          7370 => x"2e",
          7371 => x"87",
          7372 => x"76",
          7373 => x"84",
          7374 => x"80",
          7375 => x"c2",
          7376 => x"08",
          7377 => x"05",
          7378 => x"75",
          7379 => x"56",
          7380 => x"a5",
          7381 => x"fc",
          7382 => x"53",
          7383 => x"76",
          7384 => x"bf",
          7385 => x"32",
          7386 => x"05",
          7387 => x"9f",
          7388 => x"81",
          7389 => x"56",
          7390 => x"18",
          7391 => x"88",
          7392 => x"3d",
          7393 => x"3d",
          7394 => x"11",
          7395 => x"80",
          7396 => x"38",
          7397 => x"05",
          7398 => x"8c",
          7399 => x"08",
          7400 => x"3f",
          7401 => x"08",
          7402 => x"16",
          7403 => x"09",
          7404 => x"38",
          7405 => x"55",
          7406 => x"55",
          7407 => x"ec",
          7408 => x"0d",
          7409 => x"0d",
          7410 => x"cc",
          7411 => x"73",
          7412 => x"c2",
          7413 => x"0c",
          7414 => x"04",
          7415 => x"02",
          7416 => x"33",
          7417 => x"3d",
          7418 => x"54",
          7419 => x"52",
          7420 => x"a9",
          7421 => x"ff",
          7422 => x"3d",
          7423 => x"00",
          7424 => x"ff",
          7425 => x"ff",
          7426 => x"ff",
          7427 => x"00",
          7428 => x"00",
          7429 => x"00",
          7430 => x"00",
          7431 => x"00",
          7432 => x"00",
          7433 => x"00",
          7434 => x"00",
          7435 => x"00",
          7436 => x"00",
          7437 => x"00",
          7438 => x"00",
          7439 => x"00",
          7440 => x"00",
          7441 => x"00",
          7442 => x"00",
          7443 => x"00",
          7444 => x"00",
          7445 => x"00",
          7446 => x"00",
          7447 => x"00",
          7448 => x"00",
          7449 => x"00",
          7450 => x"00",
          7451 => x"00",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"00",
          7462 => x"00",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"00",
          7467 => x"00",
          7468 => x"00",
          7469 => x"00",
          7470 => x"00",
          7471 => x"00",
          7472 => x"00",
          7473 => x"00",
          7474 => x"64",
          7475 => x"74",
          7476 => x"64",
          7477 => x"74",
          7478 => x"66",
          7479 => x"74",
          7480 => x"66",
          7481 => x"64",
          7482 => x"66",
          7483 => x"63",
          7484 => x"6d",
          7485 => x"61",
          7486 => x"6d",
          7487 => x"79",
          7488 => x"6d",
          7489 => x"66",
          7490 => x"6d",
          7491 => x"70",
          7492 => x"6d",
          7493 => x"6d",
          7494 => x"6d",
          7495 => x"68",
          7496 => x"68",
          7497 => x"68",
          7498 => x"68",
          7499 => x"63",
          7500 => x"00",
          7501 => x"6a",
          7502 => x"72",
          7503 => x"61",
          7504 => x"72",
          7505 => x"74",
          7506 => x"69",
          7507 => x"00",
          7508 => x"74",
          7509 => x"00",
          7510 => x"74",
          7511 => x"69",
          7512 => x"6d",
          7513 => x"69",
          7514 => x"6b",
          7515 => x"00",
          7516 => x"65",
          7517 => x"44",
          7518 => x"20",
          7519 => x"6f",
          7520 => x"49",
          7521 => x"72",
          7522 => x"20",
          7523 => x"6f",
          7524 => x"00",
          7525 => x"44",
          7526 => x"20",
          7527 => x"20",
          7528 => x"64",
          7529 => x"00",
          7530 => x"4e",
          7531 => x"69",
          7532 => x"66",
          7533 => x"64",
          7534 => x"4e",
          7535 => x"61",
          7536 => x"66",
          7537 => x"64",
          7538 => x"49",
          7539 => x"6c",
          7540 => x"66",
          7541 => x"6e",
          7542 => x"2e",
          7543 => x"41",
          7544 => x"73",
          7545 => x"65",
          7546 => x"64",
          7547 => x"46",
          7548 => x"20",
          7549 => x"65",
          7550 => x"20",
          7551 => x"73",
          7552 => x"0a",
          7553 => x"46",
          7554 => x"20",
          7555 => x"64",
          7556 => x"69",
          7557 => x"6c",
          7558 => x"0a",
          7559 => x"53",
          7560 => x"73",
          7561 => x"69",
          7562 => x"70",
          7563 => x"65",
          7564 => x"64",
          7565 => x"44",
          7566 => x"65",
          7567 => x"6d",
          7568 => x"20",
          7569 => x"69",
          7570 => x"6c",
          7571 => x"0a",
          7572 => x"44",
          7573 => x"20",
          7574 => x"20",
          7575 => x"62",
          7576 => x"2e",
          7577 => x"4e",
          7578 => x"6f",
          7579 => x"74",
          7580 => x"65",
          7581 => x"6c",
          7582 => x"73",
          7583 => x"20",
          7584 => x"6e",
          7585 => x"6e",
          7586 => x"73",
          7587 => x"00",
          7588 => x"46",
          7589 => x"61",
          7590 => x"62",
          7591 => x"65",
          7592 => x"00",
          7593 => x"54",
          7594 => x"6f",
          7595 => x"20",
          7596 => x"72",
          7597 => x"6f",
          7598 => x"61",
          7599 => x"6c",
          7600 => x"2e",
          7601 => x"46",
          7602 => x"20",
          7603 => x"6c",
          7604 => x"65",
          7605 => x"00",
          7606 => x"49",
          7607 => x"66",
          7608 => x"69",
          7609 => x"20",
          7610 => x"6f",
          7611 => x"0a",
          7612 => x"54",
          7613 => x"6d",
          7614 => x"20",
          7615 => x"6e",
          7616 => x"6c",
          7617 => x"0a",
          7618 => x"50",
          7619 => x"6d",
          7620 => x"72",
          7621 => x"6e",
          7622 => x"72",
          7623 => x"2e",
          7624 => x"53",
          7625 => x"65",
          7626 => x"0a",
          7627 => x"55",
          7628 => x"6f",
          7629 => x"65",
          7630 => x"72",
          7631 => x"0a",
          7632 => x"20",
          7633 => x"65",
          7634 => x"73",
          7635 => x"20",
          7636 => x"20",
          7637 => x"65",
          7638 => x"65",
          7639 => x"00",
          7640 => x"72",
          7641 => x"00",
          7642 => x"25",
          7643 => x"00",
          7644 => x"3a",
          7645 => x"25",
          7646 => x"00",
          7647 => x"20",
          7648 => x"20",
          7649 => x"00",
          7650 => x"25",
          7651 => x"00",
          7652 => x"20",
          7653 => x"20",
          7654 => x"7c",
          7655 => x"7a",
          7656 => x"0a",
          7657 => x"25",
          7658 => x"00",
          7659 => x"30",
          7660 => x"35",
          7661 => x"32",
          7662 => x"76",
          7663 => x"32",
          7664 => x"20",
          7665 => x"2c",
          7666 => x"76",
          7667 => x"32",
          7668 => x"25",
          7669 => x"73",
          7670 => x"0a",
          7671 => x"5a",
          7672 => x"49",
          7673 => x"72",
          7674 => x"74",
          7675 => x"6e",
          7676 => x"72",
          7677 => x"54",
          7678 => x"72",
          7679 => x"74",
          7680 => x"75",
          7681 => x"00",
          7682 => x"50",
          7683 => x"69",
          7684 => x"72",
          7685 => x"74",
          7686 => x"49",
          7687 => x"4c",
          7688 => x"20",
          7689 => x"65",
          7690 => x"70",
          7691 => x"49",
          7692 => x"4c",
          7693 => x"20",
          7694 => x"65",
          7695 => x"70",
          7696 => x"55",
          7697 => x"30",
          7698 => x"20",
          7699 => x"65",
          7700 => x"70",
          7701 => x"55",
          7702 => x"30",
          7703 => x"20",
          7704 => x"65",
          7705 => x"70",
          7706 => x"55",
          7707 => x"31",
          7708 => x"20",
          7709 => x"65",
          7710 => x"70",
          7711 => x"55",
          7712 => x"31",
          7713 => x"20",
          7714 => x"65",
          7715 => x"70",
          7716 => x"53",
          7717 => x"69",
          7718 => x"75",
          7719 => x"69",
          7720 => x"2e",
          7721 => x"00",
          7722 => x"45",
          7723 => x"6c",
          7724 => x"20",
          7725 => x"65",
          7726 => x"2e",
          7727 => x"61",
          7728 => x"65",
          7729 => x"2e",
          7730 => x"00",
          7731 => x"7a",
          7732 => x"68",
          7733 => x"30",
          7734 => x"46",
          7735 => x"65",
          7736 => x"6f",
          7737 => x"69",
          7738 => x"6c",
          7739 => x"20",
          7740 => x"63",
          7741 => x"20",
          7742 => x"70",
          7743 => x"73",
          7744 => x"6e",
          7745 => x"6d",
          7746 => x"61",
          7747 => x"2e",
          7748 => x"2a",
          7749 => x"43",
          7750 => x"72",
          7751 => x"2e",
          7752 => x"00",
          7753 => x"43",
          7754 => x"69",
          7755 => x"2e",
          7756 => x"43",
          7757 => x"61",
          7758 => x"67",
          7759 => x"00",
          7760 => x"25",
          7761 => x"78",
          7762 => x"38",
          7763 => x"3e",
          7764 => x"6c",
          7765 => x"30",
          7766 => x"0a",
          7767 => x"44",
          7768 => x"20",
          7769 => x"6f",
          7770 => x"00",
          7771 => x"0a",
          7772 => x"70",
          7773 => x"65",
          7774 => x"25",
          7775 => x"20",
          7776 => x"58",
          7777 => x"3f",
          7778 => x"00",
          7779 => x"25",
          7780 => x"20",
          7781 => x"58",
          7782 => x"25",
          7783 => x"20",
          7784 => x"58",
          7785 => x"45",
          7786 => x"75",
          7787 => x"67",
          7788 => x"64",
          7789 => x"20",
          7790 => x"78",
          7791 => x"2e",
          7792 => x"43",
          7793 => x"69",
          7794 => x"63",
          7795 => x"20",
          7796 => x"30",
          7797 => x"2e",
          7798 => x"00",
          7799 => x"43",
          7800 => x"20",
          7801 => x"75",
          7802 => x"64",
          7803 => x"64",
          7804 => x"25",
          7805 => x"0a",
          7806 => x"52",
          7807 => x"61",
          7808 => x"6e",
          7809 => x"70",
          7810 => x"63",
          7811 => x"6f",
          7812 => x"2e",
          7813 => x"43",
          7814 => x"20",
          7815 => x"6f",
          7816 => x"6e",
          7817 => x"2e",
          7818 => x"5a",
          7819 => x"62",
          7820 => x"25",
          7821 => x"25",
          7822 => x"73",
          7823 => x"00",
          7824 => x"25",
          7825 => x"25",
          7826 => x"73",
          7827 => x"25",
          7828 => x"25",
          7829 => x"42",
          7830 => x"63",
          7831 => x"61",
          7832 => x"0a",
          7833 => x"52",
          7834 => x"69",
          7835 => x"2e",
          7836 => x"45",
          7837 => x"6c",
          7838 => x"20",
          7839 => x"65",
          7840 => x"70",
          7841 => x"2e",
          7842 => x"25",
          7843 => x"64",
          7844 => x"20",
          7845 => x"25",
          7846 => x"64",
          7847 => x"25",
          7848 => x"53",
          7849 => x"43",
          7850 => x"69",
          7851 => x"61",
          7852 => x"6e",
          7853 => x"20",
          7854 => x"6f",
          7855 => x"6f",
          7856 => x"6f",
          7857 => x"67",
          7858 => x"3a",
          7859 => x"76",
          7860 => x"73",
          7861 => x"70",
          7862 => x"65",
          7863 => x"64",
          7864 => x"20",
          7865 => x"57",
          7866 => x"44",
          7867 => x"20",
          7868 => x"30",
          7869 => x"25",
          7870 => x"29",
          7871 => x"20",
          7872 => x"53",
          7873 => x"4d",
          7874 => x"20",
          7875 => x"30",
          7876 => x"25",
          7877 => x"29",
          7878 => x"20",
          7879 => x"49",
          7880 => x"20",
          7881 => x"4d",
          7882 => x"30",
          7883 => x"25",
          7884 => x"29",
          7885 => x"20",
          7886 => x"42",
          7887 => x"20",
          7888 => x"20",
          7889 => x"30",
          7890 => x"25",
          7891 => x"29",
          7892 => x"20",
          7893 => x"52",
          7894 => x"20",
          7895 => x"20",
          7896 => x"30",
          7897 => x"25",
          7898 => x"29",
          7899 => x"20",
          7900 => x"53",
          7901 => x"41",
          7902 => x"20",
          7903 => x"65",
          7904 => x"65",
          7905 => x"25",
          7906 => x"29",
          7907 => x"20",
          7908 => x"54",
          7909 => x"52",
          7910 => x"20",
          7911 => x"69",
          7912 => x"73",
          7913 => x"25",
          7914 => x"29",
          7915 => x"20",
          7916 => x"49",
          7917 => x"20",
          7918 => x"4c",
          7919 => x"68",
          7920 => x"65",
          7921 => x"25",
          7922 => x"29",
          7923 => x"20",
          7924 => x"57",
          7925 => x"42",
          7926 => x"20",
          7927 => x"0a",
          7928 => x"20",
          7929 => x"57",
          7930 => x"32",
          7931 => x"20",
          7932 => x"49",
          7933 => x"4c",
          7934 => x"20",
          7935 => x"50",
          7936 => x"00",
          7937 => x"20",
          7938 => x"53",
          7939 => x"00",
          7940 => x"41",
          7941 => x"65",
          7942 => x"73",
          7943 => x"20",
          7944 => x"43",
          7945 => x"52",
          7946 => x"74",
          7947 => x"63",
          7948 => x"20",
          7949 => x"72",
          7950 => x"20",
          7951 => x"30",
          7952 => x"00",
          7953 => x"20",
          7954 => x"43",
          7955 => x"4d",
          7956 => x"72",
          7957 => x"74",
          7958 => x"20",
          7959 => x"72",
          7960 => x"20",
          7961 => x"30",
          7962 => x"00",
          7963 => x"20",
          7964 => x"53",
          7965 => x"6b",
          7966 => x"61",
          7967 => x"41",
          7968 => x"65",
          7969 => x"20",
          7970 => x"20",
          7971 => x"30",
          7972 => x"00",
          7973 => x"4d",
          7974 => x"3a",
          7975 => x"20",
          7976 => x"5a",
          7977 => x"49",
          7978 => x"20",
          7979 => x"20",
          7980 => x"20",
          7981 => x"20",
          7982 => x"20",
          7983 => x"30",
          7984 => x"00",
          7985 => x"20",
          7986 => x"53",
          7987 => x"65",
          7988 => x"6c",
          7989 => x"20",
          7990 => x"71",
          7991 => x"20",
          7992 => x"20",
          7993 => x"64",
          7994 => x"34",
          7995 => x"7a",
          7996 => x"20",
          7997 => x"53",
          7998 => x"4d",
          7999 => x"6f",
          8000 => x"46",
          8001 => x"20",
          8002 => x"20",
          8003 => x"20",
          8004 => x"64",
          8005 => x"34",
          8006 => x"7a",
          8007 => x"20",
          8008 => x"57",
          8009 => x"62",
          8010 => x"20",
          8011 => x"41",
          8012 => x"6c",
          8013 => x"20",
          8014 => x"71",
          8015 => x"64",
          8016 => x"34",
          8017 => x"7a",
          8018 => x"53",
          8019 => x"6c",
          8020 => x"4d",
          8021 => x"75",
          8022 => x"46",
          8023 => x"00",
          8024 => x"45",
          8025 => x"45",
          8026 => x"69",
          8027 => x"55",
          8028 => x"6f",
          8029 => x"00",
          8030 => x"01",
          8031 => x"00",
          8032 => x"00",
          8033 => x"01",
          8034 => x"00",
          8035 => x"00",
          8036 => x"01",
          8037 => x"00",
          8038 => x"00",
          8039 => x"01",
          8040 => x"00",
          8041 => x"00",
          8042 => x"01",
          8043 => x"00",
          8044 => x"00",
          8045 => x"01",
          8046 => x"00",
          8047 => x"00",
          8048 => x"01",
          8049 => x"00",
          8050 => x"00",
          8051 => x"01",
          8052 => x"00",
          8053 => x"00",
          8054 => x"01",
          8055 => x"00",
          8056 => x"00",
          8057 => x"01",
          8058 => x"00",
          8059 => x"00",
          8060 => x"01",
          8061 => x"00",
          8062 => x"00",
          8063 => x"04",
          8064 => x"00",
          8065 => x"00",
          8066 => x"04",
          8067 => x"00",
          8068 => x"00",
          8069 => x"04",
          8070 => x"00",
          8071 => x"00",
          8072 => x"03",
          8073 => x"00",
          8074 => x"00",
          8075 => x"04",
          8076 => x"00",
          8077 => x"00",
          8078 => x"04",
          8079 => x"00",
          8080 => x"00",
          8081 => x"04",
          8082 => x"00",
          8083 => x"00",
          8084 => x"03",
          8085 => x"00",
          8086 => x"00",
          8087 => x"03",
          8088 => x"00",
          8089 => x"00",
          8090 => x"03",
          8091 => x"00",
          8092 => x"00",
          8093 => x"03",
          8094 => x"00",
          8095 => x"1b",
          8096 => x"1b",
          8097 => x"1b",
          8098 => x"1b",
          8099 => x"1b",
          8100 => x"1b",
          8101 => x"1b",
          8102 => x"1b",
          8103 => x"1b",
          8104 => x"1b",
          8105 => x"1b",
          8106 => x"10",
          8107 => x"0e",
          8108 => x"0d",
          8109 => x"0b",
          8110 => x"08",
          8111 => x"06",
          8112 => x"05",
          8113 => x"04",
          8114 => x"03",
          8115 => x"02",
          8116 => x"01",
          8117 => x"68",
          8118 => x"6f",
          8119 => x"68",
          8120 => x"00",
          8121 => x"21",
          8122 => x"25",
          8123 => x"20",
          8124 => x"0a",
          8125 => x"46",
          8126 => x"65",
          8127 => x"6f",
          8128 => x"73",
          8129 => x"74",
          8130 => x"68",
          8131 => x"6f",
          8132 => x"66",
          8133 => x"20",
          8134 => x"45",
          8135 => x"0a",
          8136 => x"43",
          8137 => x"6f",
          8138 => x"70",
          8139 => x"63",
          8140 => x"74",
          8141 => x"69",
          8142 => x"72",
          8143 => x"69",
          8144 => x"20",
          8145 => x"61",
          8146 => x"6e",
          8147 => x"00",
          8148 => x"53",
          8149 => x"22",
          8150 => x"3a",
          8151 => x"3e",
          8152 => x"7c",
          8153 => x"46",
          8154 => x"46",
          8155 => x"32",
          8156 => x"eb",
          8157 => x"53",
          8158 => x"35",
          8159 => x"4e",
          8160 => x"41",
          8161 => x"20",
          8162 => x"41",
          8163 => x"20",
          8164 => x"4e",
          8165 => x"41",
          8166 => x"20",
          8167 => x"41",
          8168 => x"20",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"80",
          8174 => x"8e",
          8175 => x"45",
          8176 => x"49",
          8177 => x"90",
          8178 => x"99",
          8179 => x"59",
          8180 => x"9c",
          8181 => x"41",
          8182 => x"a5",
          8183 => x"a8",
          8184 => x"ac",
          8185 => x"b0",
          8186 => x"b4",
          8187 => x"b8",
          8188 => x"bc",
          8189 => x"c0",
          8190 => x"c4",
          8191 => x"c8",
          8192 => x"cc",
          8193 => x"d0",
          8194 => x"d4",
          8195 => x"d8",
          8196 => x"dc",
          8197 => x"e0",
          8198 => x"e4",
          8199 => x"e8",
          8200 => x"ec",
          8201 => x"f0",
          8202 => x"f4",
          8203 => x"f8",
          8204 => x"fc",
          8205 => x"2b",
          8206 => x"3d",
          8207 => x"5c",
          8208 => x"3c",
          8209 => x"7f",
          8210 => x"00",
          8211 => x"00",
          8212 => x"01",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"01",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"01",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"01",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"01",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"01",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"01",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"01",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"01",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"01",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"01",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"01",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"01",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"01",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"01",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"01",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"01",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"01",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"01",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"01",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"01",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"01",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"01",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"01",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"01",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"01",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"01",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"01",
          8333 => x"01",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"05",
          8339 => x"05",
          8340 => x"05",
          8341 => x"00",
          8342 => x"01",
          8343 => x"01",
          8344 => x"01",
          8345 => x"01",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"01",
          8372 => x"00",
          8373 => x"01",
          8374 => x"00",
          8375 => x"02",
          8376 => x"00",
          8377 => x"00",
          8378 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
