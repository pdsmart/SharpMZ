zOS_SinglePortBootBRAM.vhd