-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b83ff",
          2049 => x"f80d0b0b",
          2050 => x"0b93b904",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"9d040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b9380",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b8295",
          2210 => x"bc738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93850400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b80c3",
          2219 => x"f42d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b80c5",
          2227 => x"e02d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"95040b0b",
          2317 => x"0b8ca404",
          2318 => x"0b0b0b8c",
          2319 => x"b3040b0b",
          2320 => x"0b8cc204",
          2321 => x"0b0b0b8c",
          2322 => x"d1040b0b",
          2323 => x"0b8ce004",
          2324 => x"0b0b0b8c",
          2325 => x"f0040b0b",
          2326 => x"0b8d8004",
          2327 => x"0b0b0b8d",
          2328 => x"8f040b0b",
          2329 => x"0b8d9e04",
          2330 => x"0b0b0b8d",
          2331 => x"ad040b0b",
          2332 => x"0b8dbd04",
          2333 => x"0b0b0b8d",
          2334 => x"cd040b0b",
          2335 => x"0b8ddd04",
          2336 => x"0b0b0b8d",
          2337 => x"ed040b0b",
          2338 => x"0b8dfd04",
          2339 => x"0b0b0b8e",
          2340 => x"8d040b0b",
          2341 => x"0b8e9d04",
          2342 => x"0b0b0b8e",
          2343 => x"ad040b0b",
          2344 => x"0b8ebd04",
          2345 => x"0b0b0b8e",
          2346 => x"cd040b0b",
          2347 => x"0b8edd04",
          2348 => x"0b0b0b8e",
          2349 => x"ed040b0b",
          2350 => x"0b8efd04",
          2351 => x"0b0b0b8f",
          2352 => x"8d040b0b",
          2353 => x"0b8f9d04",
          2354 => x"0b0b0b8f",
          2355 => x"ad040b0b",
          2356 => x"0b8fbd04",
          2357 => x"0b0b0b8f",
          2358 => x"cd040b0b",
          2359 => x"0b8fdd04",
          2360 => x"0b0b0b8f",
          2361 => x"ed040b0b",
          2362 => x"0b8ffd04",
          2363 => x"0b0b0b90",
          2364 => x"8d040b0b",
          2365 => x"0b909d04",
          2366 => x"0b0b0b90",
          2367 => x"ad040b0b",
          2368 => x"0b90bd04",
          2369 => x"0b0b0b90",
          2370 => x"cd040b0b",
          2371 => x"0b90dd04",
          2372 => x"0b0b0b90",
          2373 => x"ed040b0b",
          2374 => x"0b90fd04",
          2375 => x"0b0b0b91",
          2376 => x"8d040b0b",
          2377 => x"0b919d04",
          2378 => x"0b0b0b91",
          2379 => x"ad040b0b",
          2380 => x"0b91bd04",
          2381 => x"0b0b0b91",
          2382 => x"cd040b0b",
          2383 => x"0b91dd04",
          2384 => x"0b0b0b91",
          2385 => x"ed040b0b",
          2386 => x"0b91fd04",
          2387 => x"0b0b0b92",
          2388 => x"8d040b0b",
          2389 => x"0b929d04",
          2390 => x"0b0b0b92",
          2391 => x"ad040b0b",
          2392 => x"0b92bd04",
          2393 => x"0b0b0b92",
          2394 => x"cd04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0482b6a4",
          2434 => x"0c80f4fe",
          2435 => x"2d82b6a4",
          2436 => x"0882d090",
          2437 => x"0482b6a4",
          2438 => x"0cb3b22d",
          2439 => x"82b6a408",
          2440 => x"82d09004",
          2441 => x"82b6a40c",
          2442 => x"afe32d82",
          2443 => x"b6a40882",
          2444 => x"d0900482",
          2445 => x"b6a40caf",
          2446 => x"ad2d82b6",
          2447 => x"a40882d0",
          2448 => x"900482b6",
          2449 => x"a40c94ad",
          2450 => x"2d82b6a4",
          2451 => x"0882d090",
          2452 => x"0482b6a4",
          2453 => x"0cb1c22d",
          2454 => x"82b6a408",
          2455 => x"82d09004",
          2456 => x"82b6a40c",
          2457 => x"80cfcc2d",
          2458 => x"82b6a408",
          2459 => x"82d09004",
          2460 => x"82b6a40c",
          2461 => x"80c9fb2d",
          2462 => x"82b6a408",
          2463 => x"82d09004",
          2464 => x"82b6a40c",
          2465 => x"93d82d82",
          2466 => x"b6a40882",
          2467 => x"d0900482",
          2468 => x"b6a40c96",
          2469 => x"c02d82b6",
          2470 => x"a40882d0",
          2471 => x"900482b6",
          2472 => x"a40c97cd",
          2473 => x"2d82b6a4",
          2474 => x"0882d090",
          2475 => x"0482b6a4",
          2476 => x"0c80f8a8",
          2477 => x"2d82b6a4",
          2478 => x"0882d090",
          2479 => x"0482b6a4",
          2480 => x"0c80f986",
          2481 => x"2d82b6a4",
          2482 => x"0882d090",
          2483 => x"0482b6a4",
          2484 => x"0c80f0c3",
          2485 => x"2d82b6a4",
          2486 => x"0882d090",
          2487 => x"0482b6a4",
          2488 => x"0c80f2ba",
          2489 => x"2d82b6a4",
          2490 => x"0882d090",
          2491 => x"0482b6a4",
          2492 => x"0c80f3ed",
          2493 => x"2d82b6a4",
          2494 => x"0882d090",
          2495 => x"0482b6a4",
          2496 => x"0c81d89e",
          2497 => x"2d82b6a4",
          2498 => x"0882d090",
          2499 => x"0482b6a4",
          2500 => x"0c81e58f",
          2501 => x"2d82b6a4",
          2502 => x"0882d090",
          2503 => x"0482b6a4",
          2504 => x"0c81dd83",
          2505 => x"2d82b6a4",
          2506 => x"0882d090",
          2507 => x"0482b6a4",
          2508 => x"0c81e080",
          2509 => x"2d82b6a4",
          2510 => x"0882d090",
          2511 => x"0482b6a4",
          2512 => x"0c81ea9e",
          2513 => x"2d82b6a4",
          2514 => x"0882d090",
          2515 => x"0482b6a4",
          2516 => x"0c81f2fe",
          2517 => x"2d82b6a4",
          2518 => x"0882d090",
          2519 => x"0482b6a4",
          2520 => x"0c81e3f1",
          2521 => x"2d82b6a4",
          2522 => x"0882d090",
          2523 => x"0482b6a4",
          2524 => x"0c81edbd",
          2525 => x"2d82b6a4",
          2526 => x"0882d090",
          2527 => x"0482b6a4",
          2528 => x"0c81eedc",
          2529 => x"2d82b6a4",
          2530 => x"0882d090",
          2531 => x"0482b6a4",
          2532 => x"0c81eefb",
          2533 => x"2d82b6a4",
          2534 => x"0882d090",
          2535 => x"0482b6a4",
          2536 => x"0c81f6e5",
          2537 => x"2d82b6a4",
          2538 => x"0882d090",
          2539 => x"0482b6a4",
          2540 => x"0c81f4cb",
          2541 => x"2d82b6a4",
          2542 => x"0882d090",
          2543 => x"0482b6a4",
          2544 => x"0c81f9b9",
          2545 => x"2d82b6a4",
          2546 => x"0882d090",
          2547 => x"0482b6a4",
          2548 => x"0c81efff",
          2549 => x"2d82b6a4",
          2550 => x"0882d090",
          2551 => x"0482b6a4",
          2552 => x"0c81fcb9",
          2553 => x"2d82b6a4",
          2554 => x"0882d090",
          2555 => x"0482b6a4",
          2556 => x"0c81fdba",
          2557 => x"2d82b6a4",
          2558 => x"0882d090",
          2559 => x"0482b6a4",
          2560 => x"0c81e5ef",
          2561 => x"2d82b6a4",
          2562 => x"0882d090",
          2563 => x"0482b6a4",
          2564 => x"0c81e5c8",
          2565 => x"2d82b6a4",
          2566 => x"0882d090",
          2567 => x"0482b6a4",
          2568 => x"0c81e6f3",
          2569 => x"2d82b6a4",
          2570 => x"0882d090",
          2571 => x"0482b6a4",
          2572 => x"0c81f0d6",
          2573 => x"2d82b6a4",
          2574 => x"0882d090",
          2575 => x"0482b6a4",
          2576 => x"0c81feab",
          2577 => x"2d82b6a4",
          2578 => x"0882d090",
          2579 => x"0482b6a4",
          2580 => x"0c8280b5",
          2581 => x"2d82b6a4",
          2582 => x"0882d090",
          2583 => x"0482b6a4",
          2584 => x"0c8283f7",
          2585 => x"2d82b6a4",
          2586 => x"0882d090",
          2587 => x"0482b6a4",
          2588 => x"0c81d7bd",
          2589 => x"2d82b6a4",
          2590 => x"0882d090",
          2591 => x"0482b6a4",
          2592 => x"0c8286e3",
          2593 => x"2d82b6a4",
          2594 => x"0882d090",
          2595 => x"0482b6a4",
          2596 => x"0c829598",
          2597 => x"2d82b6a4",
          2598 => x"0882d090",
          2599 => x"0482b6a4",
          2600 => x"0c829384",
          2601 => x"2d82b6a4",
          2602 => x"0882d090",
          2603 => x"0482b6a4",
          2604 => x"0c81a8f8",
          2605 => x"2d82b6a4",
          2606 => x"0882d090",
          2607 => x"0482b6a4",
          2608 => x"0c81aae2",
          2609 => x"2d82b6a4",
          2610 => x"0882d090",
          2611 => x"0482b6a4",
          2612 => x"0c81acc6",
          2613 => x"2d82b6a4",
          2614 => x"0882d090",
          2615 => x"0482b6a4",
          2616 => x"0c80f0ec",
          2617 => x"2d82b6a4",
          2618 => x"0882d090",
          2619 => x"0482b6a4",
          2620 => x"0c80f290",
          2621 => x"2d82b6a4",
          2622 => x"0882d090",
          2623 => x"0482b6a4",
          2624 => x"0c80f5f3",
          2625 => x"2d82b6a4",
          2626 => x"0882d090",
          2627 => x"0482b6a4",
          2628 => x"0c80d698",
          2629 => x"2d82b6a4",
          2630 => x"0882d090",
          2631 => x"0482b6a4",
          2632 => x"0c81a38c",
          2633 => x"2d82b6a4",
          2634 => x"0882d090",
          2635 => x"0482b6a4",
          2636 => x"0c81a3b4",
          2637 => x"2d82b6a4",
          2638 => x"0882d090",
          2639 => x"0482b6a4",
          2640 => x"0c81a7ac",
          2641 => x"2d82b6a4",
          2642 => x"0882d090",
          2643 => x"0482b6a4",
          2644 => x"0c819ff6",
          2645 => x"2d82b6a4",
          2646 => x"0882d090",
          2647 => x"043c0400",
          2648 => x"00101010",
          2649 => x"10101010",
          2650 => x"10101010",
          2651 => x"10101010",
          2652 => x"10101010",
          2653 => x"10101010",
          2654 => x"10101010",
          2655 => x"10101010",
          2656 => x"53510400",
          2657 => x"007381ff",
          2658 => x"06738306",
          2659 => x"09810583",
          2660 => x"05101010",
          2661 => x"2b0772fc",
          2662 => x"060c5151",
          2663 => x"04727280",
          2664 => x"728106ff",
          2665 => x"05097206",
          2666 => x"05711052",
          2667 => x"720a100a",
          2668 => x"5372ed38",
          2669 => x"51515351",
          2670 => x"0482b698",
          2671 => x"7082cdf4",
          2672 => x"278e3880",
          2673 => x"71708405",
          2674 => x"530c0b0b",
          2675 => x"0b93bc04",
          2676 => x"8c815180",
          2677 => x"ef860400",
          2678 => x"82b6a408",
          2679 => x"0282b6a4",
          2680 => x"0cfb3d0d",
          2681 => x"82b6a408",
          2682 => x"8c057082",
          2683 => x"b6a408fc",
          2684 => x"050c82b6",
          2685 => x"a408fc05",
          2686 => x"085482b6",
          2687 => x"a4088805",
          2688 => x"085382cd",
          2689 => x"ec085254",
          2690 => x"849a3f82",
          2691 => x"b6980870",
          2692 => x"82b6a408",
          2693 => x"f8050c82",
          2694 => x"b6a408f8",
          2695 => x"05087082",
          2696 => x"b6980c51",
          2697 => x"54873d0d",
          2698 => x"82b6a40c",
          2699 => x"0482b6a4",
          2700 => x"080282b6",
          2701 => x"a40cfb3d",
          2702 => x"0d82b6a4",
          2703 => x"08900508",
          2704 => x"85113370",
          2705 => x"81327081",
          2706 => x"06515151",
          2707 => x"52718f38",
          2708 => x"800b82b6",
          2709 => x"a4088c05",
          2710 => x"08258338",
          2711 => x"8d39800b",
          2712 => x"82b6a408",
          2713 => x"f4050c81",
          2714 => x"c43982b6",
          2715 => x"a4088c05",
          2716 => x"08ff0582",
          2717 => x"b6a4088c",
          2718 => x"050c800b",
          2719 => x"82b6a408",
          2720 => x"f8050c82",
          2721 => x"b6a40888",
          2722 => x"050882b6",
          2723 => x"a408fc05",
          2724 => x"0c82b6a4",
          2725 => x"08f80508",
          2726 => x"8a2e80f6",
          2727 => x"38800b82",
          2728 => x"b6a4088c",
          2729 => x"05082580",
          2730 => x"e93882b6",
          2731 => x"a4089005",
          2732 => x"0851a090",
          2733 => x"3f82b698",
          2734 => x"087082b6",
          2735 => x"a408f805",
          2736 => x"0c5282b6",
          2737 => x"a408f805",
          2738 => x"08ff2e09",
          2739 => x"81068d38",
          2740 => x"800b82b6",
          2741 => x"a408f405",
          2742 => x"0c80d239",
          2743 => x"82b6a408",
          2744 => x"fc050882",
          2745 => x"b6a408f8",
          2746 => x"05085353",
          2747 => x"71733482",
          2748 => x"b6a4088c",
          2749 => x"0508ff05",
          2750 => x"82b6a408",
          2751 => x"8c050c82",
          2752 => x"b6a408fc",
          2753 => x"05088105",
          2754 => x"82b6a408",
          2755 => x"fc050cff",
          2756 => x"803982b6",
          2757 => x"a408fc05",
          2758 => x"08528072",
          2759 => x"3482b6a4",
          2760 => x"08880508",
          2761 => x"7082b6a4",
          2762 => x"08f4050c",
          2763 => x"5282b6a4",
          2764 => x"08f40508",
          2765 => x"82b6980c",
          2766 => x"873d0d82",
          2767 => x"b6a40c04",
          2768 => x"82b6a408",
          2769 => x"0282b6a4",
          2770 => x"0cf43d0d",
          2771 => x"860b82b6",
          2772 => x"a408e505",
          2773 => x"3482b6a4",
          2774 => x"08880508",
          2775 => x"82b6a408",
          2776 => x"e0050cfe",
          2777 => x"0a0b82b6",
          2778 => x"a408e805",
          2779 => x"0c82b6a4",
          2780 => x"08900570",
          2781 => x"82b6a408",
          2782 => x"fc050c82",
          2783 => x"b6a408fc",
          2784 => x"05085482",
          2785 => x"b6a4088c",
          2786 => x"05085382",
          2787 => x"b6a408e0",
          2788 => x"05705351",
          2789 => x"54818d3f",
          2790 => x"82b69808",
          2791 => x"7082b6a4",
          2792 => x"08dc050c",
          2793 => x"82b6a408",
          2794 => x"ec050882",
          2795 => x"b6a40888",
          2796 => x"05080551",
          2797 => x"54807434",
          2798 => x"82b6a408",
          2799 => x"dc050870",
          2800 => x"82b6980c",
          2801 => x"548e3d0d",
          2802 => x"82b6a40c",
          2803 => x"0482b6a4",
          2804 => x"080282b6",
          2805 => x"a40cfb3d",
          2806 => x"0d82b6a4",
          2807 => x"08900570",
          2808 => x"82b6a408",
          2809 => x"fc050c82",
          2810 => x"b6a408fc",
          2811 => x"05085482",
          2812 => x"b6a4088c",
          2813 => x"05085382",
          2814 => x"b6a40888",
          2815 => x"05085254",
          2816 => x"a33f82b6",
          2817 => x"98087082",
          2818 => x"b6a408f8",
          2819 => x"050c82b6",
          2820 => x"a408f805",
          2821 => x"087082b6",
          2822 => x"980c5154",
          2823 => x"873d0d82",
          2824 => x"b6a40c04",
          2825 => x"82b6a408",
          2826 => x"0282b6a4",
          2827 => x"0ced3d0d",
          2828 => x"800b82b6",
          2829 => x"a408e405",
          2830 => x"2382b6a4",
          2831 => x"08880508",
          2832 => x"53800b8c",
          2833 => x"140c82b6",
          2834 => x"a4088805",
          2835 => x"08851133",
          2836 => x"70812a70",
          2837 => x"81327081",
          2838 => x"06515151",
          2839 => x"51537280",
          2840 => x"2e8d38ff",
          2841 => x"0b82b6a4",
          2842 => x"08e0050c",
          2843 => x"96ac3982",
          2844 => x"b6a4088c",
          2845 => x"05085372",
          2846 => x"33537282",
          2847 => x"b6a408f8",
          2848 => x"05347281",
          2849 => x"ff065372",
          2850 => x"802e95fa",
          2851 => x"3882b6a4",
          2852 => x"088c0508",
          2853 => x"810582b6",
          2854 => x"a4088c05",
          2855 => x"0c82b6a4",
          2856 => x"08e40522",
          2857 => x"70810651",
          2858 => x"5372802e",
          2859 => x"958b3882",
          2860 => x"b6a408f8",
          2861 => x"053353af",
          2862 => x"732781fc",
          2863 => x"3882b6a4",
          2864 => x"08f80533",
          2865 => x"5372b926",
          2866 => x"81ee3882",
          2867 => x"b6a408f8",
          2868 => x"05335372",
          2869 => x"b02e0981",
          2870 => x"0680c538",
          2871 => x"82b6a408",
          2872 => x"e8053370",
          2873 => x"982b7098",
          2874 => x"2c515153",
          2875 => x"72b23882",
          2876 => x"b6a408e4",
          2877 => x"05227083",
          2878 => x"2a708132",
          2879 => x"70810651",
          2880 => x"51515372",
          2881 => x"802e9938",
          2882 => x"82b6a408",
          2883 => x"e4052270",
          2884 => x"82800751",
          2885 => x"537282b6",
          2886 => x"a408e405",
          2887 => x"23fed039",
          2888 => x"82b6a408",
          2889 => x"e8053370",
          2890 => x"982b7098",
          2891 => x"2c707083",
          2892 => x"2b721173",
          2893 => x"11515151",
          2894 => x"53515553",
          2895 => x"7282b6a4",
          2896 => x"08e80534",
          2897 => x"82b6a408",
          2898 => x"e8053354",
          2899 => x"82b6a408",
          2900 => x"f8053370",
          2901 => x"15d01151",
          2902 => x"51537282",
          2903 => x"b6a408e8",
          2904 => x"053482b6",
          2905 => x"a408e805",
          2906 => x"3370982b",
          2907 => x"70982c51",
          2908 => x"51537280",
          2909 => x"258b3880",
          2910 => x"ff0b82b6",
          2911 => x"a408e805",
          2912 => x"3482b6a4",
          2913 => x"08e40522",
          2914 => x"70832a70",
          2915 => x"81065151",
          2916 => x"5372fddb",
          2917 => x"3882b6a4",
          2918 => x"08e80533",
          2919 => x"70882b70",
          2920 => x"902b7090",
          2921 => x"2c70882c",
          2922 => x"51515151",
          2923 => x"537282b6",
          2924 => x"a408ec05",
          2925 => x"23fdb839",
          2926 => x"82b6a408",
          2927 => x"e4052270",
          2928 => x"832a7081",
          2929 => x"06515153",
          2930 => x"72802e9d",
          2931 => x"3882b6a4",
          2932 => x"08e80533",
          2933 => x"70982b70",
          2934 => x"982c5151",
          2935 => x"53728a38",
          2936 => x"810b82b6",
          2937 => x"a408e805",
          2938 => x"3482b6a4",
          2939 => x"08f80533",
          2940 => x"e01182b6",
          2941 => x"a408c405",
          2942 => x"0c5382b6",
          2943 => x"a408c405",
          2944 => x"0880d826",
          2945 => x"92943882",
          2946 => x"b6a408c4",
          2947 => x"05087082",
          2948 => x"2b829788",
          2949 => x"11700851",
          2950 => x"51515372",
          2951 => x"0482b6a4",
          2952 => x"08e40522",
          2953 => x"70900751",
          2954 => x"537282b6",
          2955 => x"a408e405",
          2956 => x"2382b6a4",
          2957 => x"08e40522",
          2958 => x"70a00751",
          2959 => x"537282b6",
          2960 => x"a408e405",
          2961 => x"23fca839",
          2962 => x"82b6a408",
          2963 => x"e4052270",
          2964 => x"81800751",
          2965 => x"537282b6",
          2966 => x"a408e405",
          2967 => x"23fc9039",
          2968 => x"82b6a408",
          2969 => x"e4052270",
          2970 => x"80c00751",
          2971 => x"537282b6",
          2972 => x"a408e405",
          2973 => x"23fbf839",
          2974 => x"82b6a408",
          2975 => x"e4052270",
          2976 => x"88075153",
          2977 => x"7282b6a4",
          2978 => x"08e40523",
          2979 => x"800b82b6",
          2980 => x"a408e805",
          2981 => x"34fbd839",
          2982 => x"82b6a408",
          2983 => x"e4052270",
          2984 => x"84075153",
          2985 => x"7282b6a4",
          2986 => x"08e40523",
          2987 => x"fbc139bf",
          2988 => x"0b82b6a4",
          2989 => x"08fc0534",
          2990 => x"82b6a408",
          2991 => x"ec0522ff",
          2992 => x"11515372",
          2993 => x"82b6a408",
          2994 => x"ec052380",
          2995 => x"e30b82b6",
          2996 => x"a408f805",
          2997 => x"348da839",
          2998 => x"82b6a408",
          2999 => x"90050882",
          3000 => x"b6a40890",
          3001 => x"05088405",
          3002 => x"82b6a408",
          3003 => x"90050c70",
          3004 => x"08515372",
          3005 => x"82b6a408",
          3006 => x"fc053482",
          3007 => x"b6a408ec",
          3008 => x"0522ff11",
          3009 => x"51537282",
          3010 => x"b6a408ec",
          3011 => x"05238cef",
          3012 => x"3982b6a4",
          3013 => x"08900508",
          3014 => x"82b6a408",
          3015 => x"90050884",
          3016 => x"0582b6a4",
          3017 => x"0890050c",
          3018 => x"700882b6",
          3019 => x"a408fc05",
          3020 => x"0c82b6a4",
          3021 => x"08e40522",
          3022 => x"70832a70",
          3023 => x"81065151",
          3024 => x"51537280",
          3025 => x"2eab3882",
          3026 => x"b6a408e8",
          3027 => x"05337098",
          3028 => x"2b537298",
          3029 => x"2c5382b6",
          3030 => x"a408fc05",
          3031 => x"085253a2",
          3032 => x"d83f82b6",
          3033 => x"98085372",
          3034 => x"82b6a408",
          3035 => x"f4052399",
          3036 => x"3982b6a4",
          3037 => x"08fc0508",
          3038 => x"519d8a3f",
          3039 => x"82b69808",
          3040 => x"537282b6",
          3041 => x"a408f405",
          3042 => x"2382b6a4",
          3043 => x"08ec0522",
          3044 => x"5382b6a4",
          3045 => x"08f40522",
          3046 => x"73713154",
          3047 => x"547282b6",
          3048 => x"a408ec05",
          3049 => x"238bd839",
          3050 => x"82b6a408",
          3051 => x"90050882",
          3052 => x"b6a40890",
          3053 => x"05088405",
          3054 => x"82b6a408",
          3055 => x"90050c70",
          3056 => x"0882b6a4",
          3057 => x"08fc050c",
          3058 => x"82b6a408",
          3059 => x"e4052270",
          3060 => x"832a7081",
          3061 => x"06515151",
          3062 => x"5372802e",
          3063 => x"ab3882b6",
          3064 => x"a408e805",
          3065 => x"3370982b",
          3066 => x"5372982c",
          3067 => x"5382b6a4",
          3068 => x"08fc0508",
          3069 => x"5253a1c1",
          3070 => x"3f82b698",
          3071 => x"08537282",
          3072 => x"b6a408f4",
          3073 => x"05239939",
          3074 => x"82b6a408",
          3075 => x"fc050851",
          3076 => x"9bf33f82",
          3077 => x"b6980853",
          3078 => x"7282b6a4",
          3079 => x"08f40523",
          3080 => x"82b6a408",
          3081 => x"ec052253",
          3082 => x"82b6a408",
          3083 => x"f4052273",
          3084 => x"71315454",
          3085 => x"7282b6a4",
          3086 => x"08ec0523",
          3087 => x"8ac13982",
          3088 => x"b6a408e4",
          3089 => x"05227082",
          3090 => x"2a708106",
          3091 => x"51515372",
          3092 => x"802ea438",
          3093 => x"82b6a408",
          3094 => x"90050882",
          3095 => x"b6a40890",
          3096 => x"05088405",
          3097 => x"82b6a408",
          3098 => x"90050c70",
          3099 => x"0882b6a4",
          3100 => x"08dc050c",
          3101 => x"53a23982",
          3102 => x"b6a40890",
          3103 => x"050882b6",
          3104 => x"a4089005",
          3105 => x"08840582",
          3106 => x"b6a40890",
          3107 => x"050c7008",
          3108 => x"82b6a408",
          3109 => x"dc050c53",
          3110 => x"82b6a408",
          3111 => x"dc050882",
          3112 => x"b6a408fc",
          3113 => x"050c82b6",
          3114 => x"a408fc05",
          3115 => x"088025a4",
          3116 => x"3882b6a4",
          3117 => x"08e40522",
          3118 => x"70820751",
          3119 => x"537282b6",
          3120 => x"a408e405",
          3121 => x"2382b6a4",
          3122 => x"08fc0508",
          3123 => x"3082b6a4",
          3124 => x"08fc050c",
          3125 => x"82b6a408",
          3126 => x"e4052270",
          3127 => x"ffbf0651",
          3128 => x"537282b6",
          3129 => x"a408e405",
          3130 => x"2381af39",
          3131 => x"880b82b6",
          3132 => x"a408f405",
          3133 => x"23a93982",
          3134 => x"b6a408e4",
          3135 => x"05227080",
          3136 => x"c0075153",
          3137 => x"7282b6a4",
          3138 => x"08e40523",
          3139 => x"80f80b82",
          3140 => x"b6a408f8",
          3141 => x"0534900b",
          3142 => x"82b6a408",
          3143 => x"f4052382",
          3144 => x"b6a408e4",
          3145 => x"05227082",
          3146 => x"2a708106",
          3147 => x"51515372",
          3148 => x"802ea438",
          3149 => x"82b6a408",
          3150 => x"90050882",
          3151 => x"b6a40890",
          3152 => x"05088405",
          3153 => x"82b6a408",
          3154 => x"90050c70",
          3155 => x"0882b6a4",
          3156 => x"08d8050c",
          3157 => x"53a23982",
          3158 => x"b6a40890",
          3159 => x"050882b6",
          3160 => x"a4089005",
          3161 => x"08840582",
          3162 => x"b6a40890",
          3163 => x"050c7008",
          3164 => x"82b6a408",
          3165 => x"d8050c53",
          3166 => x"82b6a408",
          3167 => x"d8050882",
          3168 => x"b6a408fc",
          3169 => x"050c82b6",
          3170 => x"a408e405",
          3171 => x"2270cf06",
          3172 => x"51537282",
          3173 => x"b6a408e4",
          3174 => x"052382b6",
          3175 => x"a80b82b6",
          3176 => x"a408f005",
          3177 => x"0c82b6a4",
          3178 => x"08f00508",
          3179 => x"82b6a408",
          3180 => x"f4052282",
          3181 => x"b6a408fc",
          3182 => x"05087155",
          3183 => x"70545654",
          3184 => x"55a3f33f",
          3185 => x"82b69808",
          3186 => x"53727534",
          3187 => x"82b6a408",
          3188 => x"f0050882",
          3189 => x"b6a408d4",
          3190 => x"050c82b6",
          3191 => x"a408f005",
          3192 => x"08703351",
          3193 => x"53897327",
          3194 => x"a43882b6",
          3195 => x"a408f005",
          3196 => x"08537233",
          3197 => x"5482b6a4",
          3198 => x"08f80533",
          3199 => x"7015df11",
          3200 => x"51515372",
          3201 => x"82b6a408",
          3202 => x"d0053497",
          3203 => x"3982b6a4",
          3204 => x"08f00508",
          3205 => x"537233b0",
          3206 => x"11515372",
          3207 => x"82b6a408",
          3208 => x"d0053482",
          3209 => x"b6a408d4",
          3210 => x"05085382",
          3211 => x"b6a408d0",
          3212 => x"05337334",
          3213 => x"82b6a408",
          3214 => x"f0050881",
          3215 => x"0582b6a4",
          3216 => x"08f0050c",
          3217 => x"82b6a408",
          3218 => x"f4052270",
          3219 => x"5382b6a4",
          3220 => x"08fc0508",
          3221 => x"5253a2ab",
          3222 => x"3f82b698",
          3223 => x"087082b6",
          3224 => x"a408fc05",
          3225 => x"0c5382b6",
          3226 => x"a408fc05",
          3227 => x"08802e84",
          3228 => x"38feb239",
          3229 => x"82b6a408",
          3230 => x"f0050882",
          3231 => x"b6a85455",
          3232 => x"72547470",
          3233 => x"75315153",
          3234 => x"7282b6a4",
          3235 => x"08fc0534",
          3236 => x"82b6a408",
          3237 => x"e4052270",
          3238 => x"b2065153",
          3239 => x"72802e94",
          3240 => x"3882b6a4",
          3241 => x"08ec0522",
          3242 => x"ff115153",
          3243 => x"7282b6a4",
          3244 => x"08ec0523",
          3245 => x"82b6a408",
          3246 => x"e4052270",
          3247 => x"862a7081",
          3248 => x"06515153",
          3249 => x"72802e80",
          3250 => x"e73882b6",
          3251 => x"a408ec05",
          3252 => x"2270902b",
          3253 => x"82b6a408",
          3254 => x"cc050c82",
          3255 => x"b6a408cc",
          3256 => x"0508902c",
          3257 => x"82b6a408",
          3258 => x"cc050c82",
          3259 => x"b6a408f4",
          3260 => x"05225153",
          3261 => x"72902e09",
          3262 => x"81069538",
          3263 => x"82b6a408",
          3264 => x"cc0508fe",
          3265 => x"05537282",
          3266 => x"b6a408c8",
          3267 => x"05239339",
          3268 => x"82b6a408",
          3269 => x"cc0508ff",
          3270 => x"05537282",
          3271 => x"b6a408c8",
          3272 => x"052382b6",
          3273 => x"a408c805",
          3274 => x"2282b6a4",
          3275 => x"08ec0523",
          3276 => x"82b6a408",
          3277 => x"e4052270",
          3278 => x"832a7081",
          3279 => x"06515153",
          3280 => x"72802e80",
          3281 => x"d03882b6",
          3282 => x"a408e805",
          3283 => x"3370982b",
          3284 => x"70982c82",
          3285 => x"b6a408fc",
          3286 => x"05335751",
          3287 => x"51537274",
          3288 => x"24973882",
          3289 => x"b6a408e4",
          3290 => x"052270f7",
          3291 => x"06515372",
          3292 => x"82b6a408",
          3293 => x"e405239d",
          3294 => x"3982b6a4",
          3295 => x"08e80533",
          3296 => x"5382b6a4",
          3297 => x"08fc0533",
          3298 => x"73713154",
          3299 => x"547282b6",
          3300 => x"a408e805",
          3301 => x"3482b6a4",
          3302 => x"08e40522",
          3303 => x"70832a70",
          3304 => x"81065151",
          3305 => x"5372802e",
          3306 => x"b13882b6",
          3307 => x"a408e805",
          3308 => x"3370882b",
          3309 => x"70902b70",
          3310 => x"902c7088",
          3311 => x"2c515151",
          3312 => x"51537254",
          3313 => x"82b6a408",
          3314 => x"ec052270",
          3315 => x"75315153",
          3316 => x"7282b6a4",
          3317 => x"08ec0523",
          3318 => x"af3982b6",
          3319 => x"a408fc05",
          3320 => x"3370882b",
          3321 => x"70902b70",
          3322 => x"902c7088",
          3323 => x"2c515151",
          3324 => x"51537254",
          3325 => x"82b6a408",
          3326 => x"ec052270",
          3327 => x"75315153",
          3328 => x"7282b6a4",
          3329 => x"08ec0523",
          3330 => x"82b6a408",
          3331 => x"e4052270",
          3332 => x"83800651",
          3333 => x"5372b038",
          3334 => x"82b6a408",
          3335 => x"ec0522ff",
          3336 => x"11545472",
          3337 => x"82b6a408",
          3338 => x"ec052373",
          3339 => x"902b7090",
          3340 => x"2c515380",
          3341 => x"73259038",
          3342 => x"82b6a408",
          3343 => x"88050852",
          3344 => x"a0518aee",
          3345 => x"3fd23982",
          3346 => x"b6a408e4",
          3347 => x"05227081",
          3348 => x"2a708106",
          3349 => x"51515372",
          3350 => x"802e9138",
          3351 => x"82b6a408",
          3352 => x"88050852",
          3353 => x"ad518aca",
          3354 => x"3f80c739",
          3355 => x"82b6a408",
          3356 => x"e4052270",
          3357 => x"842a7081",
          3358 => x"06515153",
          3359 => x"72802e90",
          3360 => x"3882b6a4",
          3361 => x"08880508",
          3362 => x"52ab518a",
          3363 => x"a53fa339",
          3364 => x"82b6a408",
          3365 => x"e4052270",
          3366 => x"852a7081",
          3367 => x"06515153",
          3368 => x"72802e8e",
          3369 => x"3882b6a4",
          3370 => x"08880508",
          3371 => x"52a0518a",
          3372 => x"813f82b6",
          3373 => x"a408e405",
          3374 => x"2270862a",
          3375 => x"70810651",
          3376 => x"51537280",
          3377 => x"2eb13882",
          3378 => x"b6a40888",
          3379 => x"050852b0",
          3380 => x"5189df3f",
          3381 => x"82b6a408",
          3382 => x"f4052253",
          3383 => x"72902e09",
          3384 => x"81069438",
          3385 => x"82b6a408",
          3386 => x"88050852",
          3387 => x"82b6a408",
          3388 => x"f8053351",
          3389 => x"89bc3f82",
          3390 => x"b6a408e4",
          3391 => x"05227088",
          3392 => x"2a708106",
          3393 => x"51515372",
          3394 => x"802eb038",
          3395 => x"82b6a408",
          3396 => x"ec0522ff",
          3397 => x"11545472",
          3398 => x"82b6a408",
          3399 => x"ec052373",
          3400 => x"902b7090",
          3401 => x"2c515380",
          3402 => x"73259038",
          3403 => x"82b6a408",
          3404 => x"88050852",
          3405 => x"b05188fa",
          3406 => x"3fd23982",
          3407 => x"b6a408e4",
          3408 => x"05227083",
          3409 => x"2a708106",
          3410 => x"51515372",
          3411 => x"802eb038",
          3412 => x"82b6a408",
          3413 => x"e80533ff",
          3414 => x"11545472",
          3415 => x"82b6a408",
          3416 => x"e8053473",
          3417 => x"982b7098",
          3418 => x"2c515380",
          3419 => x"73259038",
          3420 => x"82b6a408",
          3421 => x"88050852",
          3422 => x"b05188b6",
          3423 => x"3fd23982",
          3424 => x"b6a408e4",
          3425 => x"05227087",
          3426 => x"2a708106",
          3427 => x"51515372",
          3428 => x"b03882b6",
          3429 => x"a408ec05",
          3430 => x"22ff1154",
          3431 => x"547282b6",
          3432 => x"a408ec05",
          3433 => x"2373902b",
          3434 => x"70902c51",
          3435 => x"53807325",
          3436 => x"903882b6",
          3437 => x"a4088805",
          3438 => x"0852a051",
          3439 => x"87f43fd2",
          3440 => x"3982b6a4",
          3441 => x"08f80533",
          3442 => x"537280e3",
          3443 => x"2e098106",
          3444 => x"973882b6",
          3445 => x"a4088805",
          3446 => x"085282b6",
          3447 => x"a408fc05",
          3448 => x"335187ce",
          3449 => x"3f81ee39",
          3450 => x"82b6a408",
          3451 => x"f8053353",
          3452 => x"7280f32e",
          3453 => x"09810680",
          3454 => x"cb3882b6",
          3455 => x"a408f405",
          3456 => x"22ff1151",
          3457 => x"537282b6",
          3458 => x"a408f405",
          3459 => x"237283ff",
          3460 => x"ff065372",
          3461 => x"83ffff2e",
          3462 => x"81bb3882",
          3463 => x"b6a40888",
          3464 => x"05085282",
          3465 => x"b6a408fc",
          3466 => x"05087033",
          3467 => x"5282b6a4",
          3468 => x"08fc0508",
          3469 => x"810582b6",
          3470 => x"a408fc05",
          3471 => x"0c5386f2",
          3472 => x"3fffb739",
          3473 => x"82b6a408",
          3474 => x"f8053353",
          3475 => x"7280d32e",
          3476 => x"09810680",
          3477 => x"cb3882b6",
          3478 => x"a408f405",
          3479 => x"22ff1151",
          3480 => x"537282b6",
          3481 => x"a408f405",
          3482 => x"237283ff",
          3483 => x"ff065372",
          3484 => x"83ffff2e",
          3485 => x"80df3882",
          3486 => x"b6a40888",
          3487 => x"05085282",
          3488 => x"b6a408fc",
          3489 => x"05087033",
          3490 => x"525386a6",
          3491 => x"3f82b6a4",
          3492 => x"08fc0508",
          3493 => x"810582b6",
          3494 => x"a408fc05",
          3495 => x"0cffb739",
          3496 => x"82b6a408",
          3497 => x"f0050882",
          3498 => x"b6a82ea9",
          3499 => x"3882b6a4",
          3500 => x"08880508",
          3501 => x"5282b6a4",
          3502 => x"08f00508",
          3503 => x"ff0582b6",
          3504 => x"a408f005",
          3505 => x"0c82b6a4",
          3506 => x"08f00508",
          3507 => x"70335253",
          3508 => x"85e03fcc",
          3509 => x"3982b6a4",
          3510 => x"08e40522",
          3511 => x"70872a70",
          3512 => x"81065151",
          3513 => x"5372802e",
          3514 => x"80c33882",
          3515 => x"b6a408ec",
          3516 => x"0522ff11",
          3517 => x"54547282",
          3518 => x"b6a408ec",
          3519 => x"05237390",
          3520 => x"2b70902c",
          3521 => x"51538073",
          3522 => x"25a33882",
          3523 => x"b6a40888",
          3524 => x"050852a0",
          3525 => x"51859b3f",
          3526 => x"d23982b6",
          3527 => x"a4088805",
          3528 => x"085282b6",
          3529 => x"a408f805",
          3530 => x"33518586",
          3531 => x"3f800b82",
          3532 => x"b6a408e4",
          3533 => x"0523eab7",
          3534 => x"3982b6a4",
          3535 => x"08f80533",
          3536 => x"5372a52e",
          3537 => x"098106a8",
          3538 => x"38810b82",
          3539 => x"b6a408e4",
          3540 => x"0523800b",
          3541 => x"82b6a408",
          3542 => x"ec052380",
          3543 => x"0b82b6a4",
          3544 => x"08e80534",
          3545 => x"8a0b82b6",
          3546 => x"a408f405",
          3547 => x"23ea8039",
          3548 => x"82b6a408",
          3549 => x"88050852",
          3550 => x"82b6a408",
          3551 => x"f8053351",
          3552 => x"84b03fe9",
          3553 => x"ea3982b6",
          3554 => x"a4088805",
          3555 => x"088c1108",
          3556 => x"7082b6a4",
          3557 => x"08e0050c",
          3558 => x"515382b6",
          3559 => x"a408e005",
          3560 => x"0882b698",
          3561 => x"0c953d0d",
          3562 => x"82b6a40c",
          3563 => x"0482b6a4",
          3564 => x"080282b6",
          3565 => x"a40cfd3d",
          3566 => x"0d82cde8",
          3567 => x"085382b6",
          3568 => x"a4088c05",
          3569 => x"085282b6",
          3570 => x"a4088805",
          3571 => x"0851e4dd",
          3572 => x"3f82b698",
          3573 => x"087082b6",
          3574 => x"980c5485",
          3575 => x"3d0d82b6",
          3576 => x"a40c0482",
          3577 => x"b6a40802",
          3578 => x"82b6a40c",
          3579 => x"fb3d0d80",
          3580 => x"0b82b6a4",
          3581 => x"08f8050c",
          3582 => x"82cdec08",
          3583 => x"85113370",
          3584 => x"812a7081",
          3585 => x"32708106",
          3586 => x"51515151",
          3587 => x"5372802e",
          3588 => x"8d38ff0b",
          3589 => x"82b6a408",
          3590 => x"f4050c81",
          3591 => x"923982b6",
          3592 => x"a4088805",
          3593 => x"08537233",
          3594 => x"82b6a408",
          3595 => x"88050881",
          3596 => x"0582b6a4",
          3597 => x"0888050c",
          3598 => x"537282b6",
          3599 => x"a408fc05",
          3600 => x"347281ff",
          3601 => x"06537280",
          3602 => x"2eb03882",
          3603 => x"cdec0882",
          3604 => x"cdec0853",
          3605 => x"82b6a408",
          3606 => x"fc053352",
          3607 => x"90110851",
          3608 => x"53722d82",
          3609 => x"b6980853",
          3610 => x"72802eff",
          3611 => x"b138ff0b",
          3612 => x"82b6a408",
          3613 => x"f8050cff",
          3614 => x"a53982cd",
          3615 => x"ec0882cd",
          3616 => x"ec085353",
          3617 => x"8a519013",
          3618 => x"0853722d",
          3619 => x"82b69808",
          3620 => x"5372802e",
          3621 => x"8a38ff0b",
          3622 => x"82b6a408",
          3623 => x"f8050c82",
          3624 => x"b6a408f8",
          3625 => x"05087082",
          3626 => x"b6a408f4",
          3627 => x"050c5382",
          3628 => x"b6a408f4",
          3629 => x"050882b6",
          3630 => x"980c873d",
          3631 => x"0d82b6a4",
          3632 => x"0c0482b6",
          3633 => x"a4080282",
          3634 => x"b6a40cfb",
          3635 => x"3d0d800b",
          3636 => x"82b6a408",
          3637 => x"f8050c82",
          3638 => x"b6a4088c",
          3639 => x"05088511",
          3640 => x"3370812a",
          3641 => x"70813270",
          3642 => x"81065151",
          3643 => x"51515372",
          3644 => x"802e8d38",
          3645 => x"ff0b82b6",
          3646 => x"a408f405",
          3647 => x"0c80f339",
          3648 => x"82b6a408",
          3649 => x"88050853",
          3650 => x"723382b6",
          3651 => x"a4088805",
          3652 => x"08810582",
          3653 => x"b6a40888",
          3654 => x"050c5372",
          3655 => x"82b6a408",
          3656 => x"fc053472",
          3657 => x"81ff0653",
          3658 => x"72802eb6",
          3659 => x"3882b6a4",
          3660 => x"088c0508",
          3661 => x"82b6a408",
          3662 => x"8c050853",
          3663 => x"82b6a408",
          3664 => x"fc053352",
          3665 => x"90110851",
          3666 => x"53722d82",
          3667 => x"b6980853",
          3668 => x"72802eff",
          3669 => x"ab38ff0b",
          3670 => x"82b6a408",
          3671 => x"f8050cff",
          3672 => x"9f3982b6",
          3673 => x"a408f805",
          3674 => x"087082b6",
          3675 => x"a408f405",
          3676 => x"0c5382b6",
          3677 => x"a408f405",
          3678 => x"0882b698",
          3679 => x"0c873d0d",
          3680 => x"82b6a40c",
          3681 => x"0482b6a4",
          3682 => x"080282b6",
          3683 => x"a40cfe3d",
          3684 => x"0d82cdec",
          3685 => x"085282b6",
          3686 => x"a4088805",
          3687 => x"0851933f",
          3688 => x"82b69808",
          3689 => x"7082b698",
          3690 => x"0c53843d",
          3691 => x"0d82b6a4",
          3692 => x"0c0482b6",
          3693 => x"a4080282",
          3694 => x"b6a40cfb",
          3695 => x"3d0d82b6",
          3696 => x"a4088c05",
          3697 => x"08851133",
          3698 => x"70812a70",
          3699 => x"81327081",
          3700 => x"06515151",
          3701 => x"51537280",
          3702 => x"2e8d38ff",
          3703 => x"0b82b6a4",
          3704 => x"08fc050c",
          3705 => x"81cb3982",
          3706 => x"b6a4088c",
          3707 => x"05088511",
          3708 => x"3370822a",
          3709 => x"70810651",
          3710 => x"51515372",
          3711 => x"802e80db",
          3712 => x"3882b6a4",
          3713 => x"088c0508",
          3714 => x"82b6a408",
          3715 => x"8c050854",
          3716 => x"548c1408",
          3717 => x"88140825",
          3718 => x"9f3882b6",
          3719 => x"a4088c05",
          3720 => x"08700870",
          3721 => x"82b6a408",
          3722 => x"88050852",
          3723 => x"57545472",
          3724 => x"75347308",
          3725 => x"8105740c",
          3726 => x"82b6a408",
          3727 => x"8c05088c",
          3728 => x"11088105",
          3729 => x"8c120c82",
          3730 => x"b6a40888",
          3731 => x"05087082",
          3732 => x"b6a408fc",
          3733 => x"050c5153",
          3734 => x"80d73982",
          3735 => x"b6a4088c",
          3736 => x"050882b6",
          3737 => x"a4088c05",
          3738 => x"085382b6",
          3739 => x"a4088805",
          3740 => x"087081ff",
          3741 => x"06539012",
          3742 => x"08515454",
          3743 => x"722d82b6",
          3744 => x"98085372",
          3745 => x"a33882b6",
          3746 => x"a4088c05",
          3747 => x"088c1108",
          3748 => x"81058c12",
          3749 => x"0c82b6a4",
          3750 => x"08880508",
          3751 => x"7082b6a4",
          3752 => x"08fc050c",
          3753 => x"51538a39",
          3754 => x"ff0b82b6",
          3755 => x"a408fc05",
          3756 => x"0c82b6a4",
          3757 => x"08fc0508",
          3758 => x"82b6980c",
          3759 => x"873d0d82",
          3760 => x"b6a40c04",
          3761 => x"82b6a408",
          3762 => x"0282b6a4",
          3763 => x"0cf93d0d",
          3764 => x"82b6a408",
          3765 => x"88050885",
          3766 => x"11337081",
          3767 => x"32708106",
          3768 => x"51515152",
          3769 => x"71802e8d",
          3770 => x"38ff0b82",
          3771 => x"b6a408f8",
          3772 => x"050c8394",
          3773 => x"3982b6a4",
          3774 => x"08880508",
          3775 => x"85113370",
          3776 => x"862a7081",
          3777 => x"06515151",
          3778 => x"5271802e",
          3779 => x"80c53882",
          3780 => x"b6a40888",
          3781 => x"050882b6",
          3782 => x"a4088805",
          3783 => x"08535385",
          3784 => x"123370ff",
          3785 => x"bf065152",
          3786 => x"71851434",
          3787 => x"82b6a408",
          3788 => x"8805088c",
          3789 => x"11088105",
          3790 => x"8c120c82",
          3791 => x"b6a40888",
          3792 => x"05088411",
          3793 => x"337082b6",
          3794 => x"a408f805",
          3795 => x"0c515152",
          3796 => x"82b63982",
          3797 => x"b6a40888",
          3798 => x"05088511",
          3799 => x"3370822a",
          3800 => x"70810651",
          3801 => x"51515271",
          3802 => x"802e80d7",
          3803 => x"3882b6a4",
          3804 => x"08880508",
          3805 => x"70087033",
          3806 => x"82b6a408",
          3807 => x"fc050c51",
          3808 => x"5282b6a4",
          3809 => x"08fc0508",
          3810 => x"a93882b6",
          3811 => x"a4088805",
          3812 => x"0882b6a4",
          3813 => x"08880508",
          3814 => x"53538512",
          3815 => x"3370a007",
          3816 => x"51527185",
          3817 => x"1434ff0b",
          3818 => x"82b6a408",
          3819 => x"f8050c81",
          3820 => x"d73982b6",
          3821 => x"a4088805",
          3822 => x"08700881",
          3823 => x"05710c52",
          3824 => x"81a13982",
          3825 => x"b6a40888",
          3826 => x"050882b6",
          3827 => x"a4088805",
          3828 => x"08529411",
          3829 => x"08515271",
          3830 => x"2d82b698",
          3831 => x"087082b6",
          3832 => x"a408fc05",
          3833 => x"0c5282b6",
          3834 => x"a408fc05",
          3835 => x"08802580",
          3836 => x"f23882b6",
          3837 => x"a4088805",
          3838 => x"0882b6a4",
          3839 => x"08f4050c",
          3840 => x"82b6a408",
          3841 => x"88050885",
          3842 => x"113382b6",
          3843 => x"a408f005",
          3844 => x"0c5282b6",
          3845 => x"a408fc05",
          3846 => x"08ff2e09",
          3847 => x"81069538",
          3848 => x"82b6a408",
          3849 => x"f0050890",
          3850 => x"07527182",
          3851 => x"b6a408ec",
          3852 => x"05349339",
          3853 => x"82b6a408",
          3854 => x"f00508a0",
          3855 => x"07527182",
          3856 => x"b6a408ec",
          3857 => x"053482b6",
          3858 => x"a408f405",
          3859 => x"085282b6",
          3860 => x"a408ec05",
          3861 => x"33851334",
          3862 => x"ff0b82b6",
          3863 => x"a408f805",
          3864 => x"0ca63982",
          3865 => x"b6a40888",
          3866 => x"05088c11",
          3867 => x"0881058c",
          3868 => x"120c82b6",
          3869 => x"a408fc05",
          3870 => x"087081ff",
          3871 => x"067082b6",
          3872 => x"a408f805",
          3873 => x"0c515152",
          3874 => x"82b6a408",
          3875 => x"f8050882",
          3876 => x"b6980c89",
          3877 => x"3d0d82b6",
          3878 => x"a40c0482",
          3879 => x"b6a40802",
          3880 => x"82b6a40c",
          3881 => x"fd3d0d82",
          3882 => x"b6a40888",
          3883 => x"050882b6",
          3884 => x"a408fc05",
          3885 => x"0c82b6a4",
          3886 => x"088c0508",
          3887 => x"82b6a408",
          3888 => x"f8050c82",
          3889 => x"b6a40890",
          3890 => x"0508802e",
          3891 => x"82a23882",
          3892 => x"b6a408f8",
          3893 => x"050882b6",
          3894 => x"a408fc05",
          3895 => x"082681ac",
          3896 => x"3882b6a4",
          3897 => x"08f80508",
          3898 => x"82b6a408",
          3899 => x"90050805",
          3900 => x"5182b6a4",
          3901 => x"08fc0508",
          3902 => x"71278190",
          3903 => x"3882b6a4",
          3904 => x"08fc0508",
          3905 => x"82b6a408",
          3906 => x"90050805",
          3907 => x"82b6a408",
          3908 => x"fc050c82",
          3909 => x"b6a408f8",
          3910 => x"050882b6",
          3911 => x"a4089005",
          3912 => x"080582b6",
          3913 => x"a408f805",
          3914 => x"0c82b6a4",
          3915 => x"08900508",
          3916 => x"810582b6",
          3917 => x"a4089005",
          3918 => x"0c82b6a4",
          3919 => x"08900508",
          3920 => x"ff0582b6",
          3921 => x"a4089005",
          3922 => x"0c82b6a4",
          3923 => x"08900508",
          3924 => x"802e819c",
          3925 => x"3882b6a4",
          3926 => x"08fc0508",
          3927 => x"ff0582b6",
          3928 => x"a408fc05",
          3929 => x"0c82b6a4",
          3930 => x"08f80508",
          3931 => x"ff0582b6",
          3932 => x"a408f805",
          3933 => x"0c82b6a4",
          3934 => x"08fc0508",
          3935 => x"82b6a408",
          3936 => x"f8050853",
          3937 => x"51713371",
          3938 => x"34ffae39",
          3939 => x"82b6a408",
          3940 => x"90050881",
          3941 => x"0582b6a4",
          3942 => x"0890050c",
          3943 => x"82b6a408",
          3944 => x"900508ff",
          3945 => x"0582b6a4",
          3946 => x"0890050c",
          3947 => x"82b6a408",
          3948 => x"90050880",
          3949 => x"2eba3882",
          3950 => x"b6a408f8",
          3951 => x"05085170",
          3952 => x"3382b6a4",
          3953 => x"08f80508",
          3954 => x"810582b6",
          3955 => x"a408f805",
          3956 => x"0c82b6a4",
          3957 => x"08fc0508",
          3958 => x"52527171",
          3959 => x"3482b6a4",
          3960 => x"08fc0508",
          3961 => x"810582b6",
          3962 => x"a408fc05",
          3963 => x"0cffad39",
          3964 => x"82b6a408",
          3965 => x"88050870",
          3966 => x"82b6980c",
          3967 => x"51853d0d",
          3968 => x"82b6a40c",
          3969 => x"0482b6a4",
          3970 => x"080282b6",
          3971 => x"a40cfe3d",
          3972 => x"0d82b6a4",
          3973 => x"08880508",
          3974 => x"82b6a408",
          3975 => x"fc050c82",
          3976 => x"b6a408fc",
          3977 => x"05085271",
          3978 => x"3382b6a4",
          3979 => x"08fc0508",
          3980 => x"810582b6",
          3981 => x"a408fc05",
          3982 => x"0c7081ff",
          3983 => x"06515170",
          3984 => x"802e8338",
          3985 => x"da3982b6",
          3986 => x"a408fc05",
          3987 => x"08ff0582",
          3988 => x"b6a408fc",
          3989 => x"050c82b6",
          3990 => x"a408fc05",
          3991 => x"0882b6a4",
          3992 => x"08880508",
          3993 => x"317082b6",
          3994 => x"980c5184",
          3995 => x"3d0d82b6",
          3996 => x"a40c0482",
          3997 => x"b6a40802",
          3998 => x"82b6a40c",
          3999 => x"fe3d0d82",
          4000 => x"b6a40888",
          4001 => x"050882b6",
          4002 => x"a408fc05",
          4003 => x"0c82b6a4",
          4004 => x"088c0508",
          4005 => x"52713382",
          4006 => x"b6a4088c",
          4007 => x"05088105",
          4008 => x"82b6a408",
          4009 => x"8c050c82",
          4010 => x"b6a408fc",
          4011 => x"05085351",
          4012 => x"70723482",
          4013 => x"b6a408fc",
          4014 => x"05088105",
          4015 => x"82b6a408",
          4016 => x"fc050c70",
          4017 => x"81ff0651",
          4018 => x"70802e84",
          4019 => x"38ffbe39",
          4020 => x"82b6a408",
          4021 => x"88050870",
          4022 => x"82b6980c",
          4023 => x"51843d0d",
          4024 => x"82b6a40c",
          4025 => x"0482b6a4",
          4026 => x"080282b6",
          4027 => x"a40cfd3d",
          4028 => x"0d82b6a4",
          4029 => x"08880508",
          4030 => x"82b6a408",
          4031 => x"fc050c82",
          4032 => x"b6a4088c",
          4033 => x"050882b6",
          4034 => x"a408f805",
          4035 => x"0c82b6a4",
          4036 => x"08900508",
          4037 => x"802e80e5",
          4038 => x"3882b6a4",
          4039 => x"08900508",
          4040 => x"810582b6",
          4041 => x"a4089005",
          4042 => x"0c82b6a4",
          4043 => x"08900508",
          4044 => x"ff0582b6",
          4045 => x"a4089005",
          4046 => x"0c82b6a4",
          4047 => x"08900508",
          4048 => x"802eba38",
          4049 => x"82b6a408",
          4050 => x"f8050851",
          4051 => x"703382b6",
          4052 => x"a408f805",
          4053 => x"08810582",
          4054 => x"b6a408f8",
          4055 => x"050c82b6",
          4056 => x"a408fc05",
          4057 => x"08525271",
          4058 => x"713482b6",
          4059 => x"a408fc05",
          4060 => x"08810582",
          4061 => x"b6a408fc",
          4062 => x"050cffad",
          4063 => x"3982b6a4",
          4064 => x"08880508",
          4065 => x"7082b698",
          4066 => x"0c51853d",
          4067 => x"0d82b6a4",
          4068 => x"0c0482b6",
          4069 => x"a4080282",
          4070 => x"b6a40cfd",
          4071 => x"3d0d82b6",
          4072 => x"a4089005",
          4073 => x"08802e81",
          4074 => x"f43882b6",
          4075 => x"a4088c05",
          4076 => x"08527133",
          4077 => x"82b6a408",
          4078 => x"8c050881",
          4079 => x"0582b6a4",
          4080 => x"088c050c",
          4081 => x"82b6a408",
          4082 => x"88050870",
          4083 => x"337281ff",
          4084 => x"06535454",
          4085 => x"5171712e",
          4086 => x"843880ce",
          4087 => x"3982b6a4",
          4088 => x"08880508",
          4089 => x"52713382",
          4090 => x"b6a40888",
          4091 => x"05088105",
          4092 => x"82b6a408",
          4093 => x"88050c70",
          4094 => x"81ff0651",
          4095 => x"51708d38",
          4096 => x"800b82b6",
          4097 => x"a408fc05",
          4098 => x"0c819b39",
          4099 => x"82b6a408",
          4100 => x"900508ff",
          4101 => x"0582b6a4",
          4102 => x"0890050c",
          4103 => x"82b6a408",
          4104 => x"90050880",
          4105 => x"2e8438ff",
          4106 => x"813982b6",
          4107 => x"a4089005",
          4108 => x"08802e80",
          4109 => x"e83882b6",
          4110 => x"a4088805",
          4111 => x"08703352",
          4112 => x"53708d38",
          4113 => x"ff0b82b6",
          4114 => x"a408fc05",
          4115 => x"0c80d739",
          4116 => x"82b6a408",
          4117 => x"8c0508ff",
          4118 => x"0582b6a4",
          4119 => x"088c050c",
          4120 => x"82b6a408",
          4121 => x"8c050870",
          4122 => x"33525270",
          4123 => x"8c38810b",
          4124 => x"82b6a408",
          4125 => x"fc050cae",
          4126 => x"3982b6a4",
          4127 => x"08880508",
          4128 => x"703382b6",
          4129 => x"a4088c05",
          4130 => x"08703372",
          4131 => x"71317082",
          4132 => x"b6a408fc",
          4133 => x"050c5355",
          4134 => x"5252538a",
          4135 => x"39800b82",
          4136 => x"b6a408fc",
          4137 => x"050c82b6",
          4138 => x"a408fc05",
          4139 => x"0882b698",
          4140 => x"0c853d0d",
          4141 => x"82b6a40c",
          4142 => x"0482b6a4",
          4143 => x"080282b6",
          4144 => x"a40cfd3d",
          4145 => x"0d82b6a4",
          4146 => x"08880508",
          4147 => x"82b6a408",
          4148 => x"f8050c82",
          4149 => x"b6a4088c",
          4150 => x"05088d38",
          4151 => x"800b82b6",
          4152 => x"a408fc05",
          4153 => x"0c80ec39",
          4154 => x"82b6a408",
          4155 => x"f8050852",
          4156 => x"713382b6",
          4157 => x"a408f805",
          4158 => x"08810582",
          4159 => x"b6a408f8",
          4160 => x"050c7081",
          4161 => x"ff065151",
          4162 => x"70802e9f",
          4163 => x"3882b6a4",
          4164 => x"088c0508",
          4165 => x"ff0582b6",
          4166 => x"a4088c05",
          4167 => x"0c82b6a4",
          4168 => x"088c0508",
          4169 => x"ff2e8438",
          4170 => x"ffbe3982",
          4171 => x"b6a408f8",
          4172 => x"0508ff05",
          4173 => x"82b6a408",
          4174 => x"f8050c82",
          4175 => x"b6a408f8",
          4176 => x"050882b6",
          4177 => x"a4088805",
          4178 => x"08317082",
          4179 => x"b6a408fc",
          4180 => x"050c5182",
          4181 => x"b6a408fc",
          4182 => x"050882b6",
          4183 => x"980c853d",
          4184 => x"0d82b6a4",
          4185 => x"0c0482b6",
          4186 => x"a4080282",
          4187 => x"b6a40cfe",
          4188 => x"3d0d82b6",
          4189 => x"a4088805",
          4190 => x"0882b6a4",
          4191 => x"08fc050c",
          4192 => x"82b6a408",
          4193 => x"90050880",
          4194 => x"2e80d438",
          4195 => x"82b6a408",
          4196 => x"90050881",
          4197 => x"0582b6a4",
          4198 => x"0890050c",
          4199 => x"82b6a408",
          4200 => x"900508ff",
          4201 => x"0582b6a4",
          4202 => x"0890050c",
          4203 => x"82b6a408",
          4204 => x"90050880",
          4205 => x"2ea93882",
          4206 => x"b6a4088c",
          4207 => x"05085170",
          4208 => x"82b6a408",
          4209 => x"fc050852",
          4210 => x"52717134",
          4211 => x"82b6a408",
          4212 => x"fc050881",
          4213 => x"0582b6a4",
          4214 => x"08fc050c",
          4215 => x"ffbe3982",
          4216 => x"b6a40888",
          4217 => x"05087082",
          4218 => x"b6980c51",
          4219 => x"843d0d82",
          4220 => x"b6a40c04",
          4221 => x"82b6a408",
          4222 => x"0282b6a4",
          4223 => x"0cf93d0d",
          4224 => x"800b82b6",
          4225 => x"a408fc05",
          4226 => x"0c82b6a4",
          4227 => x"08880508",
          4228 => x"8025b938",
          4229 => x"82b6a408",
          4230 => x"88050830",
          4231 => x"82b6a408",
          4232 => x"88050c80",
          4233 => x"0b82b6a4",
          4234 => x"08f4050c",
          4235 => x"82b6a408",
          4236 => x"fc05088a",
          4237 => x"38810b82",
          4238 => x"b6a408f4",
          4239 => x"050c82b6",
          4240 => x"a408f405",
          4241 => x"0882b6a4",
          4242 => x"08fc050c",
          4243 => x"82b6a408",
          4244 => x"8c050880",
          4245 => x"25b93882",
          4246 => x"b6a4088c",
          4247 => x"05083082",
          4248 => x"b6a4088c",
          4249 => x"050c800b",
          4250 => x"82b6a408",
          4251 => x"f0050c82",
          4252 => x"b6a408fc",
          4253 => x"05088a38",
          4254 => x"810b82b6",
          4255 => x"a408f005",
          4256 => x"0c82b6a4",
          4257 => x"08f00508",
          4258 => x"82b6a408",
          4259 => x"fc050c80",
          4260 => x"5382b6a4",
          4261 => x"088c0508",
          4262 => x"5282b6a4",
          4263 => x"08880508",
          4264 => x"5182c53f",
          4265 => x"82b69808",
          4266 => x"7082b6a4",
          4267 => x"08f8050c",
          4268 => x"5482b6a4",
          4269 => x"08fc0508",
          4270 => x"802e9038",
          4271 => x"82b6a408",
          4272 => x"f8050830",
          4273 => x"82b6a408",
          4274 => x"f8050c82",
          4275 => x"b6a408f8",
          4276 => x"05087082",
          4277 => x"b6980c54",
          4278 => x"893d0d82",
          4279 => x"b6a40c04",
          4280 => x"82b6a408",
          4281 => x"0282b6a4",
          4282 => x"0cfb3d0d",
          4283 => x"800b82b6",
          4284 => x"a408fc05",
          4285 => x"0c82b6a4",
          4286 => x"08880508",
          4287 => x"80259938",
          4288 => x"82b6a408",
          4289 => x"88050830",
          4290 => x"82b6a408",
          4291 => x"88050c81",
          4292 => x"0b82b6a4",
          4293 => x"08fc050c",
          4294 => x"82b6a408",
          4295 => x"8c050880",
          4296 => x"25903882",
          4297 => x"b6a4088c",
          4298 => x"05083082",
          4299 => x"b6a4088c",
          4300 => x"050c8153",
          4301 => x"82b6a408",
          4302 => x"8c050852",
          4303 => x"82b6a408",
          4304 => x"88050851",
          4305 => x"81a23f82",
          4306 => x"b6980870",
          4307 => x"82b6a408",
          4308 => x"f8050c54",
          4309 => x"82b6a408",
          4310 => x"fc050880",
          4311 => x"2e903882",
          4312 => x"b6a408f8",
          4313 => x"05083082",
          4314 => x"b6a408f8",
          4315 => x"050c82b6",
          4316 => x"a408f805",
          4317 => x"087082b6",
          4318 => x"980c5487",
          4319 => x"3d0d82b6",
          4320 => x"a40c0482",
          4321 => x"b6a40802",
          4322 => x"82b6a40c",
          4323 => x"fd3d0d80",
          4324 => x"5382b6a4",
          4325 => x"088c0508",
          4326 => x"5282b6a4",
          4327 => x"08880508",
          4328 => x"5180c53f",
          4329 => x"82b69808",
          4330 => x"7082b698",
          4331 => x"0c54853d",
          4332 => x"0d82b6a4",
          4333 => x"0c0482b6",
          4334 => x"a4080282",
          4335 => x"b6a40cfd",
          4336 => x"3d0d8153",
          4337 => x"82b6a408",
          4338 => x"8c050852",
          4339 => x"82b6a408",
          4340 => x"88050851",
          4341 => x"933f82b6",
          4342 => x"98087082",
          4343 => x"b6980c54",
          4344 => x"853d0d82",
          4345 => x"b6a40c04",
          4346 => x"82b6a408",
          4347 => x"0282b6a4",
          4348 => x"0cfd3d0d",
          4349 => x"810b82b6",
          4350 => x"a408fc05",
          4351 => x"0c800b82",
          4352 => x"b6a408f8",
          4353 => x"050c82b6",
          4354 => x"a4088c05",
          4355 => x"0882b6a4",
          4356 => x"08880508",
          4357 => x"27b93882",
          4358 => x"b6a408fc",
          4359 => x"0508802e",
          4360 => x"ae38800b",
          4361 => x"82b6a408",
          4362 => x"8c050824",
          4363 => x"a23882b6",
          4364 => x"a4088c05",
          4365 => x"081082b6",
          4366 => x"a4088c05",
          4367 => x"0c82b6a4",
          4368 => x"08fc0508",
          4369 => x"1082b6a4",
          4370 => x"08fc050c",
          4371 => x"ffb83982",
          4372 => x"b6a408fc",
          4373 => x"0508802e",
          4374 => x"80e13882",
          4375 => x"b6a4088c",
          4376 => x"050882b6",
          4377 => x"a4088805",
          4378 => x"0826ad38",
          4379 => x"82b6a408",
          4380 => x"88050882",
          4381 => x"b6a4088c",
          4382 => x"05083182",
          4383 => x"b6a40888",
          4384 => x"050c82b6",
          4385 => x"a408f805",
          4386 => x"0882b6a4",
          4387 => x"08fc0508",
          4388 => x"0782b6a4",
          4389 => x"08f8050c",
          4390 => x"82b6a408",
          4391 => x"fc050881",
          4392 => x"2a82b6a4",
          4393 => x"08fc050c",
          4394 => x"82b6a408",
          4395 => x"8c050881",
          4396 => x"2a82b6a4",
          4397 => x"088c050c",
          4398 => x"ff953982",
          4399 => x"b6a40890",
          4400 => x"0508802e",
          4401 => x"933882b6",
          4402 => x"a4088805",
          4403 => x"087082b6",
          4404 => x"a408f405",
          4405 => x"0c519139",
          4406 => x"82b6a408",
          4407 => x"f8050870",
          4408 => x"82b6a408",
          4409 => x"f4050c51",
          4410 => x"82b6a408",
          4411 => x"f4050882",
          4412 => x"b6980c85",
          4413 => x"3d0d82b6",
          4414 => x"a40c0482",
          4415 => x"b6a40802",
          4416 => x"82b6a40c",
          4417 => x"f73d0d80",
          4418 => x"0b82b6a4",
          4419 => x"08f00534",
          4420 => x"82b6a408",
          4421 => x"8c050853",
          4422 => x"80730c82",
          4423 => x"b6a40888",
          4424 => x"05087008",
          4425 => x"51537233",
          4426 => x"537282b6",
          4427 => x"a408f805",
          4428 => x"347281ff",
          4429 => x"065372a0",
          4430 => x"2e098106",
          4431 => x"913882b6",
          4432 => x"a4088805",
          4433 => x"08700881",
          4434 => x"05710c53",
          4435 => x"ce3982b6",
          4436 => x"a408f805",
          4437 => x"335372ad",
          4438 => x"2e098106",
          4439 => x"a438810b",
          4440 => x"82b6a408",
          4441 => x"f0053482",
          4442 => x"b6a40888",
          4443 => x"05087008",
          4444 => x"8105710c",
          4445 => x"70085153",
          4446 => x"723382b6",
          4447 => x"a408f805",
          4448 => x"3482b6a4",
          4449 => x"08f80533",
          4450 => x"5372b02e",
          4451 => x"09810681",
          4452 => x"dc3882b6",
          4453 => x"a4088805",
          4454 => x"08700881",
          4455 => x"05710c70",
          4456 => x"08515372",
          4457 => x"3382b6a4",
          4458 => x"08f80534",
          4459 => x"82b6a408",
          4460 => x"f8053382",
          4461 => x"b6a408e8",
          4462 => x"050c82b6",
          4463 => x"a408e805",
          4464 => x"0880e22e",
          4465 => x"b63882b6",
          4466 => x"a408e805",
          4467 => x"0880f82e",
          4468 => x"843880cd",
          4469 => x"39900b82",
          4470 => x"b6a408f4",
          4471 => x"053482b6",
          4472 => x"a4088805",
          4473 => x"08700881",
          4474 => x"05710c70",
          4475 => x"08515372",
          4476 => x"3382b6a4",
          4477 => x"08f80534",
          4478 => x"81a43982",
          4479 => x"0b82b6a4",
          4480 => x"08f40534",
          4481 => x"82b6a408",
          4482 => x"88050870",
          4483 => x"08810571",
          4484 => x"0c700851",
          4485 => x"53723382",
          4486 => x"b6a408f8",
          4487 => x"053480fe",
          4488 => x"3982b6a4",
          4489 => x"08f80533",
          4490 => x"5372a026",
          4491 => x"8d38810b",
          4492 => x"82b6a408",
          4493 => x"ec050c83",
          4494 => x"803982b6",
          4495 => x"a408f805",
          4496 => x"3353af73",
          4497 => x"27903882",
          4498 => x"b6a408f8",
          4499 => x"05335372",
          4500 => x"b9268338",
          4501 => x"8d39800b",
          4502 => x"82b6a408",
          4503 => x"ec050c82",
          4504 => x"d839880b",
          4505 => x"82b6a408",
          4506 => x"f40534b2",
          4507 => x"3982b6a4",
          4508 => x"08f80533",
          4509 => x"53af7327",
          4510 => x"903882b6",
          4511 => x"a408f805",
          4512 => x"335372b9",
          4513 => x"2683388d",
          4514 => x"39800b82",
          4515 => x"b6a408ec",
          4516 => x"050c82a5",
          4517 => x"398a0b82",
          4518 => x"b6a408f4",
          4519 => x"0534800b",
          4520 => x"82b6a408",
          4521 => x"fc050c82",
          4522 => x"b6a408f8",
          4523 => x"053353a0",
          4524 => x"732781cf",
          4525 => x"3882b6a4",
          4526 => x"08f80533",
          4527 => x"5380e073",
          4528 => x"27943882",
          4529 => x"b6a408f8",
          4530 => x"0533e011",
          4531 => x"51537282",
          4532 => x"b6a408f8",
          4533 => x"053482b6",
          4534 => x"a408f805",
          4535 => x"33d01151",
          4536 => x"537282b6",
          4537 => x"a408f805",
          4538 => x"3482b6a4",
          4539 => x"08f80533",
          4540 => x"53907327",
          4541 => x"ad3882b6",
          4542 => x"a408f805",
          4543 => x"33f91151",
          4544 => x"537282b6",
          4545 => x"a408f805",
          4546 => x"3482b6a4",
          4547 => x"08f80533",
          4548 => x"53728926",
          4549 => x"8d38800b",
          4550 => x"82b6a408",
          4551 => x"ec050c81",
          4552 => x"983982b6",
          4553 => x"a408f805",
          4554 => x"3382b6a4",
          4555 => x"08f40533",
          4556 => x"54547274",
          4557 => x"268d3880",
          4558 => x"0b82b6a4",
          4559 => x"08ec050c",
          4560 => x"80f73982",
          4561 => x"b6a408f4",
          4562 => x"05337082",
          4563 => x"b6a408fc",
          4564 => x"05082982",
          4565 => x"b6a408f8",
          4566 => x"05337012",
          4567 => x"82b6a408",
          4568 => x"fc050c82",
          4569 => x"b6a40888",
          4570 => x"05087008",
          4571 => x"8105710c",
          4572 => x"70085151",
          4573 => x"52555372",
          4574 => x"3382b6a4",
          4575 => x"08f80534",
          4576 => x"fea53982",
          4577 => x"b6a408f0",
          4578 => x"05335372",
          4579 => x"802e9038",
          4580 => x"82b6a408",
          4581 => x"fc050830",
          4582 => x"82b6a408",
          4583 => x"fc050c82",
          4584 => x"b6a4088c",
          4585 => x"050882b6",
          4586 => x"a408fc05",
          4587 => x"08710c53",
          4588 => x"810b82b6",
          4589 => x"a408ec05",
          4590 => x"0c82b6a4",
          4591 => x"08ec0508",
          4592 => x"82b6980c",
          4593 => x"8b3d0d82",
          4594 => x"b6a40c04",
          4595 => x"82b6a408",
          4596 => x"0282b6a4",
          4597 => x"0cf73d0d",
          4598 => x"800b82b6",
          4599 => x"a408f005",
          4600 => x"3482b6a4",
          4601 => x"088c0508",
          4602 => x"5380730c",
          4603 => x"82b6a408",
          4604 => x"88050870",
          4605 => x"08515372",
          4606 => x"33537282",
          4607 => x"b6a408f8",
          4608 => x"05347281",
          4609 => x"ff065372",
          4610 => x"a02e0981",
          4611 => x"06913882",
          4612 => x"b6a40888",
          4613 => x"05087008",
          4614 => x"8105710c",
          4615 => x"53ce3982",
          4616 => x"b6a408f8",
          4617 => x"05335372",
          4618 => x"ad2e0981",
          4619 => x"06a43881",
          4620 => x"0b82b6a4",
          4621 => x"08f00534",
          4622 => x"82b6a408",
          4623 => x"88050870",
          4624 => x"08810571",
          4625 => x"0c700851",
          4626 => x"53723382",
          4627 => x"b6a408f8",
          4628 => x"053482b6",
          4629 => x"a408f805",
          4630 => x"335372b0",
          4631 => x"2e098106",
          4632 => x"81dc3882",
          4633 => x"b6a40888",
          4634 => x"05087008",
          4635 => x"8105710c",
          4636 => x"70085153",
          4637 => x"723382b6",
          4638 => x"a408f805",
          4639 => x"3482b6a4",
          4640 => x"08f80533",
          4641 => x"82b6a408",
          4642 => x"e8050c82",
          4643 => x"b6a408e8",
          4644 => x"050880e2",
          4645 => x"2eb63882",
          4646 => x"b6a408e8",
          4647 => x"050880f8",
          4648 => x"2e843880",
          4649 => x"cd39900b",
          4650 => x"82b6a408",
          4651 => x"f4053482",
          4652 => x"b6a40888",
          4653 => x"05087008",
          4654 => x"8105710c",
          4655 => x"70085153",
          4656 => x"723382b6",
          4657 => x"a408f805",
          4658 => x"3481a439",
          4659 => x"820b82b6",
          4660 => x"a408f405",
          4661 => x"3482b6a4",
          4662 => x"08880508",
          4663 => x"70088105",
          4664 => x"710c7008",
          4665 => x"51537233",
          4666 => x"82b6a408",
          4667 => x"f8053480",
          4668 => x"fe3982b6",
          4669 => x"a408f805",
          4670 => x"335372a0",
          4671 => x"268d3881",
          4672 => x"0b82b6a4",
          4673 => x"08ec050c",
          4674 => x"83803982",
          4675 => x"b6a408f8",
          4676 => x"053353af",
          4677 => x"73279038",
          4678 => x"82b6a408",
          4679 => x"f8053353",
          4680 => x"72b92683",
          4681 => x"388d3980",
          4682 => x"0b82b6a4",
          4683 => x"08ec050c",
          4684 => x"82d83988",
          4685 => x"0b82b6a4",
          4686 => x"08f40534",
          4687 => x"b23982b6",
          4688 => x"a408f805",
          4689 => x"3353af73",
          4690 => x"27903882",
          4691 => x"b6a408f8",
          4692 => x"05335372",
          4693 => x"b9268338",
          4694 => x"8d39800b",
          4695 => x"82b6a408",
          4696 => x"ec050c82",
          4697 => x"a5398a0b",
          4698 => x"82b6a408",
          4699 => x"f4053480",
          4700 => x"0b82b6a4",
          4701 => x"08fc050c",
          4702 => x"82b6a408",
          4703 => x"f8053353",
          4704 => x"a0732781",
          4705 => x"cf3882b6",
          4706 => x"a408f805",
          4707 => x"335380e0",
          4708 => x"73279438",
          4709 => x"82b6a408",
          4710 => x"f80533e0",
          4711 => x"11515372",
          4712 => x"82b6a408",
          4713 => x"f8053482",
          4714 => x"b6a408f8",
          4715 => x"0533d011",
          4716 => x"51537282",
          4717 => x"b6a408f8",
          4718 => x"053482b6",
          4719 => x"a408f805",
          4720 => x"33539073",
          4721 => x"27ad3882",
          4722 => x"b6a408f8",
          4723 => x"0533f911",
          4724 => x"51537282",
          4725 => x"b6a408f8",
          4726 => x"053482b6",
          4727 => x"a408f805",
          4728 => x"33537289",
          4729 => x"268d3880",
          4730 => x"0b82b6a4",
          4731 => x"08ec050c",
          4732 => x"81983982",
          4733 => x"b6a408f8",
          4734 => x"053382b6",
          4735 => x"a408f405",
          4736 => x"33545472",
          4737 => x"74268d38",
          4738 => x"800b82b6",
          4739 => x"a408ec05",
          4740 => x"0c80f739",
          4741 => x"82b6a408",
          4742 => x"f4053370",
          4743 => x"82b6a408",
          4744 => x"fc050829",
          4745 => x"82b6a408",
          4746 => x"f8053370",
          4747 => x"1282b6a4",
          4748 => x"08fc050c",
          4749 => x"82b6a408",
          4750 => x"88050870",
          4751 => x"08810571",
          4752 => x"0c700851",
          4753 => x"51525553",
          4754 => x"723382b6",
          4755 => x"a408f805",
          4756 => x"34fea539",
          4757 => x"82b6a408",
          4758 => x"f0053353",
          4759 => x"72802e90",
          4760 => x"3882b6a4",
          4761 => x"08fc0508",
          4762 => x"3082b6a4",
          4763 => x"08fc050c",
          4764 => x"82b6a408",
          4765 => x"8c050882",
          4766 => x"b6a408fc",
          4767 => x"0508710c",
          4768 => x"53810b82",
          4769 => x"b6a408ec",
          4770 => x"050c82b6",
          4771 => x"a408ec05",
          4772 => x"0882b698",
          4773 => x"0c8b3d0d",
          4774 => x"82b6a40c",
          4775 => x"04f93d0d",
          4776 => x"79700870",
          4777 => x"56565874",
          4778 => x"802e80e3",
          4779 => x"38953975",
          4780 => x"0851e6d1",
          4781 => x"3f82b698",
          4782 => x"0815780c",
          4783 => x"85163354",
          4784 => x"80cd3974",
          4785 => x"335473a0",
          4786 => x"2e098106",
          4787 => x"86388115",
          4788 => x"55f13980",
          4789 => x"57769029",
          4790 => x"82b19805",
          4791 => x"70085256",
          4792 => x"e6a33f82",
          4793 => x"b6980853",
          4794 => x"74527508",
          4795 => x"51e9a33f",
          4796 => x"82b69808",
          4797 => x"8b388416",
          4798 => x"33547381",
          4799 => x"2effb038",
          4800 => x"81177081",
          4801 => x"ff065854",
          4802 => x"997727c9",
          4803 => x"38ff5473",
          4804 => x"82b6980c",
          4805 => x"893d0d04",
          4806 => x"ff3d0d73",
          4807 => x"52719326",
          4808 => x"818e3871",
          4809 => x"84298295",
          4810 => x"cc055271",
          4811 => x"0804829b",
          4812 => x"98518180",
          4813 => x"39829ba4",
          4814 => x"5180f939",
          4815 => x"829bb451",
          4816 => x"80f23982",
          4817 => x"9bc45180",
          4818 => x"eb39829b",
          4819 => x"d45180e4",
          4820 => x"39829be4",
          4821 => x"5180dd39",
          4822 => x"829bf851",
          4823 => x"80d63982",
          4824 => x"9c885180",
          4825 => x"cf39829c",
          4826 => x"a05180c8",
          4827 => x"39829cb8",
          4828 => x"5180c139",
          4829 => x"829cd051",
          4830 => x"bb39829c",
          4831 => x"ec51b539",
          4832 => x"829d8051",
          4833 => x"af39829d",
          4834 => x"a851a939",
          4835 => x"829db851",
          4836 => x"a339829d",
          4837 => x"d8519d39",
          4838 => x"829de851",
          4839 => x"9739829e",
          4840 => x"80519139",
          4841 => x"829e9851",
          4842 => x"8b39829e",
          4843 => x"b0518539",
          4844 => x"829ebc51",
          4845 => x"d8ad3f83",
          4846 => x"3d0d04fb",
          4847 => x"3d0d7779",
          4848 => x"56567487",
          4849 => x"e7268a38",
          4850 => x"74527587",
          4851 => x"e8295190",
          4852 => x"3987e852",
          4853 => x"7451efab",
          4854 => x"3f82b698",
          4855 => x"08527551",
          4856 => x"efa13f82",
          4857 => x"b6980854",
          4858 => x"79537552",
          4859 => x"829ecc51",
          4860 => x"ffbbe53f",
          4861 => x"873d0d04",
          4862 => x"ec3d0d66",
          4863 => x"02840580",
          4864 => x"e305335b",
          4865 => x"57806878",
          4866 => x"30707a07",
          4867 => x"73255157",
          4868 => x"59597856",
          4869 => x"7787ff26",
          4870 => x"83388156",
          4871 => x"74760770",
          4872 => x"81ff0651",
          4873 => x"55935674",
          4874 => x"81823881",
          4875 => x"5376528c",
          4876 => x"3d705256",
          4877 => x"80ffe73f",
          4878 => x"82b69808",
          4879 => x"5782b698",
          4880 => x"08b93882",
          4881 => x"b6980887",
          4882 => x"c098880c",
          4883 => x"82b69808",
          4884 => x"59963dd4",
          4885 => x"05548480",
          4886 => x"53775275",
          4887 => x"518184a3",
          4888 => x"3f82b698",
          4889 => x"085782b6",
          4890 => x"98089038",
          4891 => x"7a557480",
          4892 => x"2e893874",
          4893 => x"19751959",
          4894 => x"59d73996",
          4895 => x"3dd80551",
          4896 => x"818c8c3f",
          4897 => x"76307078",
          4898 => x"0780257b",
          4899 => x"30709f2a",
          4900 => x"72065157",
          4901 => x"51567480",
          4902 => x"2e903882",
          4903 => x"9ef05387",
          4904 => x"c0988808",
          4905 => x"527851fe",
          4906 => x"923f7656",
          4907 => x"7582b698",
          4908 => x"0c963d0d",
          4909 => x"04f73d0d",
          4910 => x"7d028405",
          4911 => x"bb053359",
          4912 => x"5aff5980",
          4913 => x"537c527b",
          4914 => x"51fead3f",
          4915 => x"82b69808",
          4916 => x"80cb3877",
          4917 => x"802e8838",
          4918 => x"77812ebf",
          4919 => x"38bf3982",
          4920 => x"cde85782",
          4921 => x"cde85682",
          4922 => x"cde85582",
          4923 => x"cdf00854",
          4924 => x"82cdec08",
          4925 => x"5382cde8",
          4926 => x"0852829e",
          4927 => x"f851ffb9",
          4928 => x"d73f82cd",
          4929 => x"e8566255",
          4930 => x"615482b6",
          4931 => x"98536052",
          4932 => x"7f51792d",
          4933 => x"82b69808",
          4934 => x"59833979",
          4935 => x"047882b6",
          4936 => x"980c8b3d",
          4937 => x"0d04f33d",
          4938 => x"0d7f6163",
          4939 => x"028c0580",
          4940 => x"cf053373",
          4941 => x"73156841",
          4942 => x"5f5c5c5e",
          4943 => x"5e5e7a52",
          4944 => x"829fac51",
          4945 => x"ffb9913f",
          4946 => x"829fb451",
          4947 => x"ffb9893f",
          4948 => x"80557479",
          4949 => x"27818038",
          4950 => x"7b902e89",
          4951 => x"387ba02e",
          4952 => x"a73880c6",
          4953 => x"39741853",
          4954 => x"727a278e",
          4955 => x"38722252",
          4956 => x"829fb851",
          4957 => x"ffb8e13f",
          4958 => x"8939829f",
          4959 => x"c451ffb8",
          4960 => x"d73f8215",
          4961 => x"5580c339",
          4962 => x"74185372",
          4963 => x"7a278e38",
          4964 => x"72085282",
          4965 => x"9fac51ff",
          4966 => x"b8be3f89",
          4967 => x"39829fc0",
          4968 => x"51ffb8b4",
          4969 => x"3f841555",
          4970 => x"a1397418",
          4971 => x"53727a27",
          4972 => x"8e387233",
          4973 => x"52829fcc",
          4974 => x"51ffb89c",
          4975 => x"3f893982",
          4976 => x"9fd451ff",
          4977 => x"b8923f81",
          4978 => x"155582cd",
          4979 => x"ec0852a0",
          4980 => x"51d7df3f",
          4981 => x"fefc3982",
          4982 => x"9fd851ff",
          4983 => x"b7fa3f80",
          4984 => x"55747927",
          4985 => x"80c63874",
          4986 => x"18703355",
          4987 => x"53805672",
          4988 => x"7a278338",
          4989 => x"81568053",
          4990 => x"9f742783",
          4991 => x"38815375",
          4992 => x"73067081",
          4993 => x"ff065153",
          4994 => x"72802e90",
          4995 => x"387380fe",
          4996 => x"268a3882",
          4997 => x"cdec0852",
          4998 => x"73518839",
          4999 => x"82cdec08",
          5000 => x"52a051d7",
          5001 => x"8d3f8115",
          5002 => x"55ffb639",
          5003 => x"829fdc51",
          5004 => x"d3b13f78",
          5005 => x"18791c5c",
          5006 => x"589ccb3f",
          5007 => x"82b69808",
          5008 => x"982b7098",
          5009 => x"2c515776",
          5010 => x"a02e0981",
          5011 => x"06aa389c",
          5012 => x"b53f82b6",
          5013 => x"9808982b",
          5014 => x"70982c70",
          5015 => x"a0327030",
          5016 => x"729b3270",
          5017 => x"30707207",
          5018 => x"73750706",
          5019 => x"51585859",
          5020 => x"57515780",
          5021 => x"7324d838",
          5022 => x"769b2e09",
          5023 => x"81068538",
          5024 => x"80538c39",
          5025 => x"7c1e5372",
          5026 => x"7826fdb2",
          5027 => x"38ff5372",
          5028 => x"82b6980c",
          5029 => x"8f3d0d04",
          5030 => x"fc3d0d02",
          5031 => x"9b053382",
          5032 => x"9fe05382",
          5033 => x"9fe45255",
          5034 => x"ffb6ad3f",
          5035 => x"82b4f022",
          5036 => x"51a5a43f",
          5037 => x"829ff054",
          5038 => x"829ffc53",
          5039 => x"82b4f133",
          5040 => x"5282a084",
          5041 => x"51ffb690",
          5042 => x"3f74802e",
          5043 => x"8438a0d8",
          5044 => x"3f863d0d",
          5045 => x"04fe3d0d",
          5046 => x"87c09680",
          5047 => x"0853a5c0",
          5048 => x"3f815198",
          5049 => x"8e3f82a0",
          5050 => x"a05199a3",
          5051 => x"3f805198",
          5052 => x"823f7281",
          5053 => x"2a708106",
          5054 => x"51527180",
          5055 => x"2e923881",
          5056 => x"5197f03f",
          5057 => x"82a0b851",
          5058 => x"99853f80",
          5059 => x"5197e43f",
          5060 => x"72822a70",
          5061 => x"81065152",
          5062 => x"71802e92",
          5063 => x"38815197",
          5064 => x"d23f82a0",
          5065 => x"c85198e7",
          5066 => x"3f805197",
          5067 => x"c63f7283",
          5068 => x"2a708106",
          5069 => x"51527180",
          5070 => x"2e923881",
          5071 => x"5197b43f",
          5072 => x"82a0d851",
          5073 => x"98c93f80",
          5074 => x"5197a83f",
          5075 => x"72842a70",
          5076 => x"81065152",
          5077 => x"71802e92",
          5078 => x"38815197",
          5079 => x"963f82a0",
          5080 => x"ec5198ab",
          5081 => x"3f805197",
          5082 => x"8a3f7285",
          5083 => x"2a708106",
          5084 => x"51527180",
          5085 => x"2e923881",
          5086 => x"5196f83f",
          5087 => x"82a18051",
          5088 => x"988d3f80",
          5089 => x"5196ec3f",
          5090 => x"72862a70",
          5091 => x"81065152",
          5092 => x"71802e92",
          5093 => x"38815196",
          5094 => x"da3f82a1",
          5095 => x"945197ef",
          5096 => x"3f805196",
          5097 => x"ce3f7287",
          5098 => x"2a708106",
          5099 => x"51527180",
          5100 => x"2e923881",
          5101 => x"5196bc3f",
          5102 => x"82a1a851",
          5103 => x"97d13f80",
          5104 => x"5196b03f",
          5105 => x"72882a70",
          5106 => x"81065152",
          5107 => x"71802e92",
          5108 => x"38815196",
          5109 => x"9e3f82a1",
          5110 => x"bc5197b3",
          5111 => x"3f805196",
          5112 => x"923fa3c4",
          5113 => x"3f843d0d",
          5114 => x"04fb3d0d",
          5115 => x"77028405",
          5116 => x"a3053370",
          5117 => x"55565680",
          5118 => x"527551e2",
          5119 => x"e93f0b0b",
          5120 => x"82b19433",
          5121 => x"5473a938",
          5122 => x"815382a1",
          5123 => x"f85282cd",
          5124 => x"985180f8",
          5125 => x"893f82b6",
          5126 => x"98083070",
          5127 => x"82b69808",
          5128 => x"07802582",
          5129 => x"71315151",
          5130 => x"54730b0b",
          5131 => x"82b19434",
          5132 => x"0b0b82b1",
          5133 => x"94335473",
          5134 => x"812e0981",
          5135 => x"06af3882",
          5136 => x"cd985374",
          5137 => x"52755181",
          5138 => x"b2ba3f82",
          5139 => x"b6980880",
          5140 => x"2e8b3882",
          5141 => x"b6980851",
          5142 => x"cf893f91",
          5143 => x"3982cd98",
          5144 => x"518184ab",
          5145 => x"3f820b0b",
          5146 => x"0b82b194",
          5147 => x"340b0b82",
          5148 => x"b1943354",
          5149 => x"73822e09",
          5150 => x"81068c38",
          5151 => x"82a28853",
          5152 => x"74527551",
          5153 => x"a9bc3f80",
          5154 => x"0b82b698",
          5155 => x"0c873d0d",
          5156 => x"04ce3d0d",
          5157 => x"80707182",
          5158 => x"cd940c5f",
          5159 => x"5d81527c",
          5160 => x"5180c6d5",
          5161 => x"3f82b698",
          5162 => x"0881ff06",
          5163 => x"59787d2e",
          5164 => x"098106a3",
          5165 => x"38963d59",
          5166 => x"835382a2",
          5167 => x"90527851",
          5168 => x"dca33f7c",
          5169 => x"53785282",
          5170 => x"b7c45180",
          5171 => x"f5ef3f82",
          5172 => x"b698087d",
          5173 => x"2e883882",
          5174 => x"a294518d",
          5175 => x"a3398170",
          5176 => x"5f5d82a2",
          5177 => x"cc51ffb1",
          5178 => x"ef3f963d",
          5179 => x"70465a80",
          5180 => x"f8527951",
          5181 => x"fdf33fb4",
          5182 => x"3dff8405",
          5183 => x"51f39e3f",
          5184 => x"82b69808",
          5185 => x"902b7090",
          5186 => x"2c515978",
          5187 => x"80c22e87",
          5188 => x"a3387880",
          5189 => x"c224b238",
          5190 => x"78bd2e81",
          5191 => x"d23878bd",
          5192 => x"24903878",
          5193 => x"802effba",
          5194 => x"3878bc2e",
          5195 => x"80da388a",
          5196 => x"d4397880",
          5197 => x"c02e8399",
          5198 => x"387880c0",
          5199 => x"2485cd38",
          5200 => x"78bf2e82",
          5201 => x"8c388abd",
          5202 => x"397880f9",
          5203 => x"2e89d938",
          5204 => x"7880f924",
          5205 => x"92387880",
          5206 => x"c32e8888",
          5207 => x"387880f8",
          5208 => x"2e89a138",
          5209 => x"8a9f3978",
          5210 => x"81832e8a",
          5211 => x"86387881",
          5212 => x"83248b38",
          5213 => x"7881822e",
          5214 => x"89eb388a",
          5215 => x"88397881",
          5216 => x"852e89fb",
          5217 => x"3889fe39",
          5218 => x"b43dff80",
          5219 => x"1153ff84",
          5220 => x"0551ecb8",
          5221 => x"3f82b698",
          5222 => x"08802efe",
          5223 => x"c538b43d",
          5224 => x"fefc1153",
          5225 => x"ff840551",
          5226 => x"eca23f82",
          5227 => x"b6980880",
          5228 => x"2efeaf38",
          5229 => x"b43dfef8",
          5230 => x"1153ff84",
          5231 => x"0551ec8c",
          5232 => x"3f82b698",
          5233 => x"08863882",
          5234 => x"b6980842",
          5235 => x"82a2d051",
          5236 => x"ffb0853f",
          5237 => x"63635c5a",
          5238 => x"797b2781",
          5239 => x"ec386159",
          5240 => x"787a7084",
          5241 => x"055c0c7a",
          5242 => x"7a26f538",
          5243 => x"81db39b4",
          5244 => x"3dff8011",
          5245 => x"53ff8405",
          5246 => x"51ebd13f",
          5247 => x"82b69808",
          5248 => x"802efdde",
          5249 => x"38b43dfe",
          5250 => x"fc1153ff",
          5251 => x"840551eb",
          5252 => x"bb3f82b6",
          5253 => x"9808802e",
          5254 => x"fdc838b4",
          5255 => x"3dfef811",
          5256 => x"53ff8405",
          5257 => x"51eba53f",
          5258 => x"82b69808",
          5259 => x"802efdb2",
          5260 => x"3882a2e0",
          5261 => x"51ffafa0",
          5262 => x"3f635a79",
          5263 => x"63278189",
          5264 => x"38615979",
          5265 => x"7081055b",
          5266 => x"33793461",
          5267 => x"810542eb",
          5268 => x"39b43dff",
          5269 => x"801153ff",
          5270 => x"840551ea",
          5271 => x"ef3f82b6",
          5272 => x"9808802e",
          5273 => x"fcfc38b4",
          5274 => x"3dfefc11",
          5275 => x"53ff8405",
          5276 => x"51ead93f",
          5277 => x"82b69808",
          5278 => x"802efce6",
          5279 => x"38b43dfe",
          5280 => x"f81153ff",
          5281 => x"840551ea",
          5282 => x"c33f82b6",
          5283 => x"9808802e",
          5284 => x"fcd03882",
          5285 => x"a2ec51ff",
          5286 => x"aebe3f63",
          5287 => x"5a796327",
          5288 => x"a8386170",
          5289 => x"337b335e",
          5290 => x"5a5b787c",
          5291 => x"2e923878",
          5292 => x"557a5479",
          5293 => x"33537952",
          5294 => x"82a2fc51",
          5295 => x"ffae993f",
          5296 => x"811a6281",
          5297 => x"05435ad5",
          5298 => x"398a51cd",
          5299 => x"b83ffc92",
          5300 => x"39b43dff",
          5301 => x"801153ff",
          5302 => x"840551e9",
          5303 => x"ef3f82b6",
          5304 => x"980880df",
          5305 => x"3882b584",
          5306 => x"33597880",
          5307 => x"2e893882",
          5308 => x"b4bc0844",
          5309 => x"80cd3982",
          5310 => x"b5853359",
          5311 => x"78802e88",
          5312 => x"3882b4c4",
          5313 => x"0844bc39",
          5314 => x"82b58633",
          5315 => x"5978802e",
          5316 => x"883882b4",
          5317 => x"cc0844ab",
          5318 => x"3982b587",
          5319 => x"33597880",
          5320 => x"2e883882",
          5321 => x"b4d40844",
          5322 => x"9a3982b5",
          5323 => x"82335978",
          5324 => x"802e8838",
          5325 => x"82b4dc08",
          5326 => x"44893982",
          5327 => x"b4ec08fc",
          5328 => x"800544b4",
          5329 => x"3dfefc11",
          5330 => x"53ff8405",
          5331 => x"51e8fd3f",
          5332 => x"82b69808",
          5333 => x"80de3882",
          5334 => x"b5843359",
          5335 => x"78802e89",
          5336 => x"3882b4c0",
          5337 => x"084380cc",
          5338 => x"3982b585",
          5339 => x"33597880",
          5340 => x"2e883882",
          5341 => x"b4c80843",
          5342 => x"bb3982b5",
          5343 => x"86335978",
          5344 => x"802e8838",
          5345 => x"82b4d008",
          5346 => x"43aa3982",
          5347 => x"b5873359",
          5348 => x"78802e88",
          5349 => x"3882b4d8",
          5350 => x"08439939",
          5351 => x"82b58233",
          5352 => x"5978802e",
          5353 => x"883882b4",
          5354 => x"e0084388",
          5355 => x"3982b4ec",
          5356 => x"08880543",
          5357 => x"b43dfef8",
          5358 => x"1153ff84",
          5359 => x"0551e88c",
          5360 => x"3f82b698",
          5361 => x"08802ea7",
          5362 => x"3880625c",
          5363 => x"5c7a882e",
          5364 => x"8338815c",
          5365 => x"7a903270",
          5366 => x"30707207",
          5367 => x"9f2a707f",
          5368 => x"0651515a",
          5369 => x"5a78802e",
          5370 => x"88387aa0",
          5371 => x"2e833888",
          5372 => x"4282a398",
          5373 => x"51c7ec3f",
          5374 => x"a0556354",
          5375 => x"61536252",
          5376 => x"6351f2a2",
          5377 => x"3f82a3a4",
          5378 => x"5186f539",
          5379 => x"b43dff80",
          5380 => x"1153ff84",
          5381 => x"0551e7b4",
          5382 => x"3f82b698",
          5383 => x"08802ef9",
          5384 => x"c138b43d",
          5385 => x"fefc1153",
          5386 => x"ff840551",
          5387 => x"e79e3f82",
          5388 => x"b6980880",
          5389 => x"2ea43863",
          5390 => x"590280cb",
          5391 => x"05337934",
          5392 => x"63810544",
          5393 => x"b43dfefc",
          5394 => x"1153ff84",
          5395 => x"0551e6fc",
          5396 => x"3f82b698",
          5397 => x"08e138f9",
          5398 => x"89396370",
          5399 => x"33545282",
          5400 => x"a3b051ff",
          5401 => x"aaf23f82",
          5402 => x"cde80853",
          5403 => x"80f85279",
          5404 => x"51ffabb9",
          5405 => x"3f794579",
          5406 => x"335978ae",
          5407 => x"2ef8e338",
          5408 => x"9f79279f",
          5409 => x"38b43dfe",
          5410 => x"fc1153ff",
          5411 => x"840551e6",
          5412 => x"bb3f82b6",
          5413 => x"9808802e",
          5414 => x"91386359",
          5415 => x"0280cb05",
          5416 => x"33793463",
          5417 => x"810544ff",
          5418 => x"b13982a3",
          5419 => x"bc51c6b3",
          5420 => x"3fffa739",
          5421 => x"b43dfef4",
          5422 => x"1153ff84",
          5423 => x"0551e0bb",
          5424 => x"3f82b698",
          5425 => x"08802ef8",
          5426 => x"9938b43d",
          5427 => x"fef01153",
          5428 => x"ff840551",
          5429 => x"e0a53f82",
          5430 => x"b6980880",
          5431 => x"2ea53860",
          5432 => x"5902be05",
          5433 => x"22797082",
          5434 => x"055b2378",
          5435 => x"41b43dfe",
          5436 => x"f01153ff",
          5437 => x"840551e0",
          5438 => x"823f82b6",
          5439 => x"9808e038",
          5440 => x"f7e03960",
          5441 => x"70225452",
          5442 => x"82a3c051",
          5443 => x"ffa9c93f",
          5444 => x"82cde808",
          5445 => x"5380f852",
          5446 => x"7951ffaa",
          5447 => x"903f7945",
          5448 => x"79335978",
          5449 => x"ae2ef7ba",
          5450 => x"38789f26",
          5451 => x"87386082",
          5452 => x"0541d039",
          5453 => x"b43dfef0",
          5454 => x"1153ff84",
          5455 => x"0551dfbb",
          5456 => x"3f82b698",
          5457 => x"08802e92",
          5458 => x"38605902",
          5459 => x"be052279",
          5460 => x"7082055b",
          5461 => x"237841ff",
          5462 => x"aa3982a3",
          5463 => x"bc51c583",
          5464 => x"3fffa039",
          5465 => x"b43dfef4",
          5466 => x"1153ff84",
          5467 => x"0551df8b",
          5468 => x"3f82b698",
          5469 => x"08802ef6",
          5470 => x"e938b43d",
          5471 => x"fef01153",
          5472 => x"ff840551",
          5473 => x"def53f82",
          5474 => x"b6980880",
          5475 => x"2ea03860",
          5476 => x"60710c59",
          5477 => x"60840541",
          5478 => x"b43dfef0",
          5479 => x"1153ff84",
          5480 => x"0551ded7",
          5481 => x"3f82b698",
          5482 => x"08e538f6",
          5483 => x"b5396070",
          5484 => x"08545282",
          5485 => x"a3cc51ff",
          5486 => x"a89e3f82",
          5487 => x"cde80853",
          5488 => x"80f85279",
          5489 => x"51ffa8e5",
          5490 => x"3f794579",
          5491 => x"335978ae",
          5492 => x"2ef68f38",
          5493 => x"9f79279b",
          5494 => x"38b43dfe",
          5495 => x"f01153ff",
          5496 => x"840551de",
          5497 => x"963f82b6",
          5498 => x"9808802e",
          5499 => x"8d386060",
          5500 => x"710c5960",
          5501 => x"840541ff",
          5502 => x"b53982a3",
          5503 => x"bc51c3e3",
          5504 => x"3fffab39",
          5505 => x"b43dff80",
          5506 => x"1153ff84",
          5507 => x"0551e3bc",
          5508 => x"3f82b698",
          5509 => x"08802ef5",
          5510 => x"c9386352",
          5511 => x"82a3dc51",
          5512 => x"ffa7b53f",
          5513 => x"63597804",
          5514 => x"b43dff80",
          5515 => x"1153ff84",
          5516 => x"0551e398",
          5517 => x"3f82b698",
          5518 => x"08802ef5",
          5519 => x"a5386352",
          5520 => x"82a3f851",
          5521 => x"ffa7913f",
          5522 => x"6359782d",
          5523 => x"82b69808",
          5524 => x"802ef58e",
          5525 => x"3882b698",
          5526 => x"085282a4",
          5527 => x"9451ffa6",
          5528 => x"f73ff4fe",
          5529 => x"3982a4b0",
          5530 => x"51c2f83f",
          5531 => x"ffa6ca3f",
          5532 => x"f4f03982",
          5533 => x"a4cc51c2",
          5534 => x"ea3f8059",
          5535 => x"ffa83991",
          5536 => x"a73ff4de",
          5537 => x"39794579",
          5538 => x"33597880",
          5539 => x"2ef4d338",
          5540 => x"7d7d0659",
          5541 => x"78802e81",
          5542 => x"cf38b43d",
          5543 => x"ff840551",
          5544 => x"83ca3f82",
          5545 => x"b698085c",
          5546 => x"815b7a82",
          5547 => x"2eb2387a",
          5548 => x"82248938",
          5549 => x"7a812e8c",
          5550 => x"3880ca39",
          5551 => x"7a832ead",
          5552 => x"3880c239",
          5553 => x"82a4e056",
          5554 => x"7b5582a4",
          5555 => x"e4548053",
          5556 => x"82a4e852",
          5557 => x"b43dffb0",
          5558 => x"0551ffa8",
          5559 => x"e33fb839",
          5560 => x"7b52b43d",
          5561 => x"ffb00551",
          5562 => x"cf893fab",
          5563 => x"397b5582",
          5564 => x"a4e45480",
          5565 => x"5382a4f8",
          5566 => x"52b43dff",
          5567 => x"b00551ff",
          5568 => x"a8be3f93",
          5569 => x"397b5480",
          5570 => x"5382a584",
          5571 => x"52b43dff",
          5572 => x"b00551ff",
          5573 => x"a8aa3f82",
          5574 => x"b4bc5882",
          5575 => x"b6c85780",
          5576 => x"56645580",
          5577 => x"5482d080",
          5578 => x"5382d080",
          5579 => x"52b43dff",
          5580 => x"b00551eb",
          5581 => x"803f82b6",
          5582 => x"980882b6",
          5583 => x"98080970",
          5584 => x"30707207",
          5585 => x"8025515b",
          5586 => x"5b5f805a",
          5587 => x"7a832683",
          5588 => x"38815a78",
          5589 => x"7a065978",
          5590 => x"802e8d38",
          5591 => x"811b7081",
          5592 => x"ff065c59",
          5593 => x"7afec338",
          5594 => x"7d81327d",
          5595 => x"81320759",
          5596 => x"788a387e",
          5597 => x"ff2e0981",
          5598 => x"06f2e738",
          5599 => x"82a58c51",
          5600 => x"c0e13ff2",
          5601 => x"dd39f53d",
          5602 => x"0d800b82",
          5603 => x"b6c83487",
          5604 => x"c0948c70",
          5605 => x"08545587",
          5606 => x"84805272",
          5607 => x"51d7e43f",
          5608 => x"82b69808",
          5609 => x"902b7508",
          5610 => x"55538784",
          5611 => x"80527351",
          5612 => x"d7d13f72",
          5613 => x"82b69808",
          5614 => x"07750c87",
          5615 => x"c0949c70",
          5616 => x"08545587",
          5617 => x"84805272",
          5618 => x"51d7b83f",
          5619 => x"82b69808",
          5620 => x"902b7508",
          5621 => x"55538784",
          5622 => x"80527351",
          5623 => x"d7a53f72",
          5624 => x"82b69808",
          5625 => x"07750c8c",
          5626 => x"80830b87",
          5627 => x"c094840c",
          5628 => x"8c80830b",
          5629 => x"87c09494",
          5630 => x"0c80f68b",
          5631 => x"5a80f8f7",
          5632 => x"5b830284",
          5633 => x"05990534",
          5634 => x"805c82cd",
          5635 => x"e80b873d",
          5636 => x"7088130c",
          5637 => x"70720c82",
          5638 => x"cdec0c54",
          5639 => x"89be3f92",
          5640 => x"ff3f82a5",
          5641 => x"9c51ffbf",
          5642 => x"ba3f82a5",
          5643 => x"a851ffbf",
          5644 => x"b23f80dd",
          5645 => x"d55192e3",
          5646 => x"3f8151ec",
          5647 => x"db3ff0d1",
          5648 => x"3f8004fe",
          5649 => x"3d0d8052",
          5650 => x"83537188",
          5651 => x"2b5287d8",
          5652 => x"3f82b698",
          5653 => x"0881ff06",
          5654 => x"7207ff14",
          5655 => x"54527280",
          5656 => x"25e83871",
          5657 => x"82b6980c",
          5658 => x"843d0d04",
          5659 => x"fc3d0d76",
          5660 => x"70085455",
          5661 => x"80735254",
          5662 => x"72742e81",
          5663 => x"8a387233",
          5664 => x"5170a02e",
          5665 => x"09810686",
          5666 => x"38811353",
          5667 => x"f1397233",
          5668 => x"5170a22e",
          5669 => x"09810686",
          5670 => x"38811353",
          5671 => x"81547252",
          5672 => x"73812e09",
          5673 => x"81069f38",
          5674 => x"84398112",
          5675 => x"52807233",
          5676 => x"525470a2",
          5677 => x"2e833881",
          5678 => x"5470802e",
          5679 => x"9d3873ea",
          5680 => x"38983981",
          5681 => x"12528072",
          5682 => x"33525470",
          5683 => x"a02e8338",
          5684 => x"81547080",
          5685 => x"2e843873",
          5686 => x"ea388072",
          5687 => x"33525470",
          5688 => x"a02e0981",
          5689 => x"06833881",
          5690 => x"5470a232",
          5691 => x"70307080",
          5692 => x"25760751",
          5693 => x"51517080",
          5694 => x"2e883880",
          5695 => x"72708105",
          5696 => x"54347175",
          5697 => x"0c725170",
          5698 => x"82b6980c",
          5699 => x"863d0d04",
          5700 => x"fc3d0d76",
          5701 => x"53720880",
          5702 => x"2e913886",
          5703 => x"3dfc0552",
          5704 => x"7251d7d7",
          5705 => x"3f82b698",
          5706 => x"08853880",
          5707 => x"53833974",
          5708 => x"537282b6",
          5709 => x"980c863d",
          5710 => x"0d04fc3d",
          5711 => x"0d768211",
          5712 => x"33ff0552",
          5713 => x"53815270",
          5714 => x"8b268198",
          5715 => x"38831333",
          5716 => x"ff055182",
          5717 => x"52709e26",
          5718 => x"818a3884",
          5719 => x"13335183",
          5720 => x"52709726",
          5721 => x"80fe3885",
          5722 => x"13335184",
          5723 => x"5270bb26",
          5724 => x"80f23886",
          5725 => x"13335185",
          5726 => x"5270bb26",
          5727 => x"80e63888",
          5728 => x"13225586",
          5729 => x"527487e7",
          5730 => x"2680d938",
          5731 => x"8a132254",
          5732 => x"87527387",
          5733 => x"e72680cc",
          5734 => x"38810b87",
          5735 => x"c0989c0c",
          5736 => x"722287c0",
          5737 => x"98bc0c82",
          5738 => x"133387c0",
          5739 => x"98b80c83",
          5740 => x"133387c0",
          5741 => x"98b40c84",
          5742 => x"133387c0",
          5743 => x"98b00c85",
          5744 => x"133387c0",
          5745 => x"98ac0c86",
          5746 => x"133387c0",
          5747 => x"98a80c74",
          5748 => x"87c098a4",
          5749 => x"0c7387c0",
          5750 => x"98a00c80",
          5751 => x"0b87c098",
          5752 => x"9c0c8052",
          5753 => x"7182b698",
          5754 => x"0c863d0d",
          5755 => x"04f33d0d",
          5756 => x"7f5b87c0",
          5757 => x"989c5d81",
          5758 => x"7d0c87c0",
          5759 => x"98bc085e",
          5760 => x"7d7b2387",
          5761 => x"c098b808",
          5762 => x"5a79821c",
          5763 => x"3487c098",
          5764 => x"b4085a79",
          5765 => x"831c3487",
          5766 => x"c098b008",
          5767 => x"5a79841c",
          5768 => x"3487c098",
          5769 => x"ac085a79",
          5770 => x"851c3487",
          5771 => x"c098a808",
          5772 => x"5a79861c",
          5773 => x"3487c098",
          5774 => x"a4085c7b",
          5775 => x"881c2387",
          5776 => x"c098a008",
          5777 => x"5a798a1c",
          5778 => x"23807d0c",
          5779 => x"7983ffff",
          5780 => x"06597b83",
          5781 => x"ffff0658",
          5782 => x"861b3357",
          5783 => x"851b3356",
          5784 => x"841b3355",
          5785 => x"831b3354",
          5786 => x"821b3353",
          5787 => x"7d83ffff",
          5788 => x"065282a5",
          5789 => x"c051ff9e",
          5790 => x"df3f8f3d",
          5791 => x"0d04fb3d",
          5792 => x"0d029f05",
          5793 => x"3382b4b8",
          5794 => x"337081ff",
          5795 => x"06585555",
          5796 => x"87c09484",
          5797 => x"5175802e",
          5798 => x"863887c0",
          5799 => x"94945170",
          5800 => x"0870962a",
          5801 => x"70810653",
          5802 => x"54527080",
          5803 => x"2e8c3871",
          5804 => x"912a7081",
          5805 => x"06515170",
          5806 => x"d7387281",
          5807 => x"32708106",
          5808 => x"51517080",
          5809 => x"2e8d3871",
          5810 => x"932a7081",
          5811 => x"06515170",
          5812 => x"ffbe3873",
          5813 => x"81ff0651",
          5814 => x"87c09480",
          5815 => x"5270802e",
          5816 => x"863887c0",
          5817 => x"94905274",
          5818 => x"720c7482",
          5819 => x"b6980c87",
          5820 => x"3d0d04ff",
          5821 => x"3d0d028f",
          5822 => x"05337030",
          5823 => x"709f2a51",
          5824 => x"52527082",
          5825 => x"b4b83483",
          5826 => x"3d0d04f9",
          5827 => x"3d0d02a7",
          5828 => x"05335877",
          5829 => x"8a2e0981",
          5830 => x"0687387a",
          5831 => x"528d51eb",
          5832 => x"3f82b4b8",
          5833 => x"337081ff",
          5834 => x"06585687",
          5835 => x"c0948453",
          5836 => x"76802e86",
          5837 => x"3887c094",
          5838 => x"94537208",
          5839 => x"70962a70",
          5840 => x"81065556",
          5841 => x"5472802e",
          5842 => x"8c387391",
          5843 => x"2a708106",
          5844 => x"515372d7",
          5845 => x"38748132",
          5846 => x"70810651",
          5847 => x"5372802e",
          5848 => x"8d387393",
          5849 => x"2a708106",
          5850 => x"515372ff",
          5851 => x"be387581",
          5852 => x"ff065387",
          5853 => x"c0948054",
          5854 => x"72802e86",
          5855 => x"3887c094",
          5856 => x"90547774",
          5857 => x"0c800b82",
          5858 => x"b6980c89",
          5859 => x"3d0d04f9",
          5860 => x"3d0d7954",
          5861 => x"80743370",
          5862 => x"81ff0653",
          5863 => x"53577077",
          5864 => x"2e80fc38",
          5865 => x"7181ff06",
          5866 => x"811582b4",
          5867 => x"b8337081",
          5868 => x"ff065957",
          5869 => x"555887c0",
          5870 => x"94845175",
          5871 => x"802e8638",
          5872 => x"87c09494",
          5873 => x"51700870",
          5874 => x"962a7081",
          5875 => x"06535452",
          5876 => x"70802e8c",
          5877 => x"3871912a",
          5878 => x"70810651",
          5879 => x"5170d738",
          5880 => x"72813270",
          5881 => x"81065151",
          5882 => x"70802e8d",
          5883 => x"3871932a",
          5884 => x"70810651",
          5885 => x"5170ffbe",
          5886 => x"387481ff",
          5887 => x"065187c0",
          5888 => x"94805270",
          5889 => x"802e8638",
          5890 => x"87c09490",
          5891 => x"5277720c",
          5892 => x"81177433",
          5893 => x"7081ff06",
          5894 => x"53535770",
          5895 => x"ff863876",
          5896 => x"82b6980c",
          5897 => x"893d0d04",
          5898 => x"fe3d0d82",
          5899 => x"b4b83370",
          5900 => x"81ff0654",
          5901 => x"5287c094",
          5902 => x"84517280",
          5903 => x"2e863887",
          5904 => x"c0949451",
          5905 => x"70087082",
          5906 => x"2a708106",
          5907 => x"51515170",
          5908 => x"802ee238",
          5909 => x"7181ff06",
          5910 => x"5187c094",
          5911 => x"80527080",
          5912 => x"2e863887",
          5913 => x"c0949052",
          5914 => x"71087081",
          5915 => x"ff0682b6",
          5916 => x"980c5184",
          5917 => x"3d0d04ff",
          5918 => x"af3f82b6",
          5919 => x"980881ff",
          5920 => x"0682b698",
          5921 => x"0c04fe3d",
          5922 => x"0d82b4b8",
          5923 => x"337081ff",
          5924 => x"06525387",
          5925 => x"c0948452",
          5926 => x"70802e86",
          5927 => x"3887c094",
          5928 => x"94527108",
          5929 => x"70822a70",
          5930 => x"81065151",
          5931 => x"51ff5270",
          5932 => x"802ea038",
          5933 => x"7281ff06",
          5934 => x"5187c094",
          5935 => x"80527080",
          5936 => x"2e863887",
          5937 => x"c0949052",
          5938 => x"71087098",
          5939 => x"2b70982c",
          5940 => x"51535171",
          5941 => x"82b6980c",
          5942 => x"843d0d04",
          5943 => x"ff3d0d87",
          5944 => x"c09e8008",
          5945 => x"709c2a8a",
          5946 => x"06515170",
          5947 => x"802e84b4",
          5948 => x"3887c09e",
          5949 => x"a40882b4",
          5950 => x"bc0c87c0",
          5951 => x"9ea80882",
          5952 => x"b4c00c87",
          5953 => x"c09e9408",
          5954 => x"82b4c40c",
          5955 => x"87c09e98",
          5956 => x"0882b4c8",
          5957 => x"0c87c09e",
          5958 => x"9c0882b4",
          5959 => x"cc0c87c0",
          5960 => x"9ea00882",
          5961 => x"b4d00c87",
          5962 => x"c09eac08",
          5963 => x"82b4d40c",
          5964 => x"87c09eb0",
          5965 => x"0882b4d8",
          5966 => x"0c87c09e",
          5967 => x"b40882b4",
          5968 => x"dc0c87c0",
          5969 => x"9eb80882",
          5970 => x"b4e00c87",
          5971 => x"c09ebc08",
          5972 => x"82b4e40c",
          5973 => x"87c09ec0",
          5974 => x"0882b4e8",
          5975 => x"0c87c09e",
          5976 => x"c40882b4",
          5977 => x"ec0c87c0",
          5978 => x"9e800851",
          5979 => x"7082b4f0",
          5980 => x"2387c09e",
          5981 => x"840882b4",
          5982 => x"f40c87c0",
          5983 => x"9e880882",
          5984 => x"b4f80c87",
          5985 => x"c09e8c08",
          5986 => x"82b4fc0c",
          5987 => x"810b82b5",
          5988 => x"8034800b",
          5989 => x"87c09e90",
          5990 => x"08708480",
          5991 => x"0a065152",
          5992 => x"5270802e",
          5993 => x"83388152",
          5994 => x"7182b581",
          5995 => x"34800b87",
          5996 => x"c09e9008",
          5997 => x"7088800a",
          5998 => x"06515252",
          5999 => x"70802e83",
          6000 => x"38815271",
          6001 => x"82b58234",
          6002 => x"800b87c0",
          6003 => x"9e900870",
          6004 => x"90800a06",
          6005 => x"51525270",
          6006 => x"802e8338",
          6007 => x"81527182",
          6008 => x"b5833480",
          6009 => x"0b87c09e",
          6010 => x"90087088",
          6011 => x"80800651",
          6012 => x"52527080",
          6013 => x"2e833881",
          6014 => x"527182b5",
          6015 => x"8434800b",
          6016 => x"87c09e90",
          6017 => x"0870a080",
          6018 => x"80065152",
          6019 => x"5270802e",
          6020 => x"83388152",
          6021 => x"7182b585",
          6022 => x"34800b87",
          6023 => x"c09e9008",
          6024 => x"70908080",
          6025 => x"06515252",
          6026 => x"70802e83",
          6027 => x"38815271",
          6028 => x"82b58634",
          6029 => x"800b87c0",
          6030 => x"9e900870",
          6031 => x"84808006",
          6032 => x"51525270",
          6033 => x"802e8338",
          6034 => x"81527182",
          6035 => x"b5873480",
          6036 => x"0b87c09e",
          6037 => x"90087082",
          6038 => x"80800651",
          6039 => x"52527080",
          6040 => x"2e833881",
          6041 => x"527182b5",
          6042 => x"8834800b",
          6043 => x"87c09e90",
          6044 => x"08708180",
          6045 => x"80065152",
          6046 => x"5270802e",
          6047 => x"83388152",
          6048 => x"7182b589",
          6049 => x"34800b87",
          6050 => x"c09e9008",
          6051 => x"7080c080",
          6052 => x"06515252",
          6053 => x"70802e83",
          6054 => x"38815271",
          6055 => x"82b58a34",
          6056 => x"800b87c0",
          6057 => x"9e900870",
          6058 => x"a0800651",
          6059 => x"52527080",
          6060 => x"2e833881",
          6061 => x"527182b5",
          6062 => x"8b3487c0",
          6063 => x"9e900870",
          6064 => x"98800670",
          6065 => x"8a2a5151",
          6066 => x"517082b5",
          6067 => x"8c34800b",
          6068 => x"87c09e90",
          6069 => x"08708480",
          6070 => x"06515252",
          6071 => x"70802e83",
          6072 => x"38815271",
          6073 => x"82b58d34",
          6074 => x"87c09e90",
          6075 => x"087083f0",
          6076 => x"0670842a",
          6077 => x"51515170",
          6078 => x"82b58e34",
          6079 => x"800b87c0",
          6080 => x"9e900870",
          6081 => x"88065152",
          6082 => x"5270802e",
          6083 => x"83388152",
          6084 => x"7182b58f",
          6085 => x"3487c09e",
          6086 => x"90087087",
          6087 => x"06515170",
          6088 => x"82b59034",
          6089 => x"833d0d04",
          6090 => x"fb3d0d82",
          6091 => x"a5d851ff",
          6092 => x"95a63f82",
          6093 => x"b5803354",
          6094 => x"73802e89",
          6095 => x"3882a5ec",
          6096 => x"51ff9594",
          6097 => x"3f82a680",
          6098 => x"51ffb197",
          6099 => x"3f82b582",
          6100 => x"33547380",
          6101 => x"2e943882",
          6102 => x"b4dc0882",
          6103 => x"b4e00811",
          6104 => x"545282a6",
          6105 => x"9851ff94",
          6106 => x"ef3f82b5",
          6107 => x"87335473",
          6108 => x"802e9438",
          6109 => x"82b4d408",
          6110 => x"82b4d808",
          6111 => x"11545282",
          6112 => x"a6b451ff",
          6113 => x"94d23f82",
          6114 => x"b5843354",
          6115 => x"73802e94",
          6116 => x"3882b4bc",
          6117 => x"0882b4c0",
          6118 => x"08115452",
          6119 => x"82a6d051",
          6120 => x"ff94b53f",
          6121 => x"82b58533",
          6122 => x"5473802e",
          6123 => x"943882b4",
          6124 => x"c40882b4",
          6125 => x"c8081154",
          6126 => x"5282a6ec",
          6127 => x"51ff9498",
          6128 => x"3f82b586",
          6129 => x"33547380",
          6130 => x"2e943882",
          6131 => x"b4cc0882",
          6132 => x"b4d00811",
          6133 => x"545282a7",
          6134 => x"8851ff93",
          6135 => x"fb3f82b5",
          6136 => x"8b335473",
          6137 => x"802e8e38",
          6138 => x"82b58c33",
          6139 => x"5282a7a4",
          6140 => x"51ff93e4",
          6141 => x"3f82b58f",
          6142 => x"33547380",
          6143 => x"2e8e3882",
          6144 => x"b5903352",
          6145 => x"82a7c451",
          6146 => x"ff93cd3f",
          6147 => x"82b58d33",
          6148 => x"5473802e",
          6149 => x"8e3882b5",
          6150 => x"8e335282",
          6151 => x"a7e451ff",
          6152 => x"93b63f82",
          6153 => x"b5813354",
          6154 => x"73802e89",
          6155 => x"3882a884",
          6156 => x"51ffafaf",
          6157 => x"3f82b583",
          6158 => x"33547380",
          6159 => x"2e893882",
          6160 => x"a89851ff",
          6161 => x"af9d3f82",
          6162 => x"b5883354",
          6163 => x"73802e89",
          6164 => x"3882a8a4",
          6165 => x"51ffaf8b",
          6166 => x"3f82b589",
          6167 => x"33547380",
          6168 => x"2e893882",
          6169 => x"a8b051ff",
          6170 => x"aef93f82",
          6171 => x"b58a3354",
          6172 => x"73802e89",
          6173 => x"3882a8b8",
          6174 => x"51ffaee7",
          6175 => x"3f82a8c0",
          6176 => x"51ffaedf",
          6177 => x"3f82b4e4",
          6178 => x"085282a8",
          6179 => x"cc51ff92",
          6180 => x"c73f82b4",
          6181 => x"e8085282",
          6182 => x"a8f451ff",
          6183 => x"92ba3f82",
          6184 => x"b4ec0852",
          6185 => x"82a99c51",
          6186 => x"ff92ad3f",
          6187 => x"82a9c451",
          6188 => x"ffaeb03f",
          6189 => x"82b4f022",
          6190 => x"5282a9cc",
          6191 => x"51ff9298",
          6192 => x"3f82b4f4",
          6193 => x"0856bd84",
          6194 => x"c0527551",
          6195 => x"c5b53f82",
          6196 => x"b69808bd",
          6197 => x"84c02976",
          6198 => x"71315454",
          6199 => x"82b69808",
          6200 => x"5282a9f4",
          6201 => x"51ff91f0",
          6202 => x"3f82b587",
          6203 => x"33547380",
          6204 => x"2ea93882",
          6205 => x"b4f80856",
          6206 => x"bd84c052",
          6207 => x"7551c583",
          6208 => x"3f82b698",
          6209 => x"08bd84c0",
          6210 => x"29767131",
          6211 => x"545482b6",
          6212 => x"98085282",
          6213 => x"aaa051ff",
          6214 => x"91be3f82",
          6215 => x"b5823354",
          6216 => x"73802ea9",
          6217 => x"3882b4fc",
          6218 => x"0856bd84",
          6219 => x"c0527551",
          6220 => x"c4d13f82",
          6221 => x"b69808bd",
          6222 => x"84c02976",
          6223 => x"71315454",
          6224 => x"82b69808",
          6225 => x"5282aacc",
          6226 => x"51ff918c",
          6227 => x"3f8a51ff",
          6228 => x"b0b33f87",
          6229 => x"3d0d04fe",
          6230 => x"3d0d0292",
          6231 => x"0533ff05",
          6232 => x"52718426",
          6233 => x"aa387184",
          6234 => x"2982969c",
          6235 => x"05527108",
          6236 => x"0482aaf8",
          6237 => x"519d3982",
          6238 => x"ab805197",
          6239 => x"3982ab88",
          6240 => x"51913982",
          6241 => x"ab90518b",
          6242 => x"3982ab94",
          6243 => x"51853982",
          6244 => x"ab9c51ff",
          6245 => x"90c23f84",
          6246 => x"3d0d0471",
          6247 => x"88800c04",
          6248 => x"800b87c0",
          6249 => x"96840c04",
          6250 => x"82b59408",
          6251 => x"87c09684",
          6252 => x"0c04fd3d",
          6253 => x"0d76982b",
          6254 => x"70982c79",
          6255 => x"982b7098",
          6256 => x"2c721013",
          6257 => x"70822b51",
          6258 => x"53515451",
          6259 => x"51800b82",
          6260 => x"aba81233",
          6261 => x"55537174",
          6262 => x"259c3882",
          6263 => x"aba41108",
          6264 => x"12028405",
          6265 => x"97053371",
          6266 => x"33525252",
          6267 => x"70722e09",
          6268 => x"81068338",
          6269 => x"81537282",
          6270 => x"b6980c85",
          6271 => x"3d0d04fb",
          6272 => x"3d0d7902",
          6273 => x"8405a305",
          6274 => x"33713355",
          6275 => x"56547280",
          6276 => x"2eb13882",
          6277 => x"cdec0852",
          6278 => x"8851ffaf",
          6279 => x"953f82cd",
          6280 => x"ec0852a0",
          6281 => x"51ffaf8a",
          6282 => x"3f82cdec",
          6283 => x"08528851",
          6284 => x"ffaeff3f",
          6285 => x"7333ff05",
          6286 => x"53727434",
          6287 => x"7281ff06",
          6288 => x"53cc3977",
          6289 => x"51ff8f90",
          6290 => x"3f747434",
          6291 => x"873d0d04",
          6292 => x"f63d0d7c",
          6293 => x"028405b7",
          6294 => x"05330288",
          6295 => x"05bb0533",
          6296 => x"82b5f033",
          6297 => x"70842982",
          6298 => x"b5980570",
          6299 => x"08515959",
          6300 => x"5a585974",
          6301 => x"802e8638",
          6302 => x"74519afa",
          6303 => x"3f82b5f0",
          6304 => x"33708429",
          6305 => x"82b59805",
          6306 => x"81197054",
          6307 => x"58565a9d",
          6308 => x"fb3f82b6",
          6309 => x"9808750c",
          6310 => x"82b5f033",
          6311 => x"70842982",
          6312 => x"b5980570",
          6313 => x"0851565a",
          6314 => x"74802ea7",
          6315 => x"38755378",
          6316 => x"527451ff",
          6317 => x"b8af3f82",
          6318 => x"b5f03381",
          6319 => x"05557482",
          6320 => x"b5f03474",
          6321 => x"81ff0655",
          6322 => x"93752787",
          6323 => x"38800b82",
          6324 => x"b5f03477",
          6325 => x"802eb638",
          6326 => x"82b5ec08",
          6327 => x"5675802e",
          6328 => x"ac3882b5",
          6329 => x"e8335574",
          6330 => x"a4388c3d",
          6331 => x"fc055476",
          6332 => x"53785275",
          6333 => x"5180da88",
          6334 => x"3f82b5ec",
          6335 => x"08528a51",
          6336 => x"818f953f",
          6337 => x"82b5ec08",
          6338 => x"5180dde5",
          6339 => x"3f8c3d0d",
          6340 => x"04fd3d0d",
          6341 => x"82b59853",
          6342 => x"93547208",
          6343 => x"5271802e",
          6344 => x"89387151",
          6345 => x"99d03f80",
          6346 => x"730cff14",
          6347 => x"84145454",
          6348 => x"738025e6",
          6349 => x"38800b82",
          6350 => x"b5f03482",
          6351 => x"b5ec0852",
          6352 => x"71802e95",
          6353 => x"38715180",
          6354 => x"dec53f82",
          6355 => x"b5ec0851",
          6356 => x"99a43f80",
          6357 => x"0b82b5ec",
          6358 => x"0c853d0d",
          6359 => x"04dc3d0d",
          6360 => x"81578052",
          6361 => x"82b5ec08",
          6362 => x"5180e3b2",
          6363 => x"3f82b698",
          6364 => x"0880d338",
          6365 => x"82b5ec08",
          6366 => x"5380f852",
          6367 => x"883d7052",
          6368 => x"56818c80",
          6369 => x"3f82b698",
          6370 => x"08802eba",
          6371 => x"387551ff",
          6372 => x"b4f33f82",
          6373 => x"b6980855",
          6374 => x"800b82b6",
          6375 => x"9808259d",
          6376 => x"3882b698",
          6377 => x"08ff0570",
          6378 => x"17555580",
          6379 => x"74347553",
          6380 => x"76528117",
          6381 => x"82ae9852",
          6382 => x"57ff8c9c",
          6383 => x"3f74ff2e",
          6384 => x"098106ff",
          6385 => x"af38a63d",
          6386 => x"0d04d93d",
          6387 => x"0daa3d08",
          6388 => x"ad3d085a",
          6389 => x"5a817058",
          6390 => x"58805282",
          6391 => x"b5ec0851",
          6392 => x"80e2bb3f",
          6393 => x"82b69808",
          6394 => x"819538ff",
          6395 => x"0b82b5ec",
          6396 => x"08545580",
          6397 => x"f8528b3d",
          6398 => x"70525681",
          6399 => x"8b863f82",
          6400 => x"b6980880",
          6401 => x"2ea53875",
          6402 => x"51ffb3f9",
          6403 => x"3f82b698",
          6404 => x"08811858",
          6405 => x"55800b82",
          6406 => x"b6980825",
          6407 => x"8e3882b6",
          6408 => x"9808ff05",
          6409 => x"70175555",
          6410 => x"80743474",
          6411 => x"09703070",
          6412 => x"72079f2a",
          6413 => x"51555578",
          6414 => x"772e8538",
          6415 => x"73ffac38",
          6416 => x"82b5ec08",
          6417 => x"8c110853",
          6418 => x"5180e1d2",
          6419 => x"3f82b698",
          6420 => x"08802e89",
          6421 => x"3882aea4",
          6422 => x"51ff8afc",
          6423 => x"3f78772e",
          6424 => x"0981069b",
          6425 => x"38755279",
          6426 => x"51ffb487",
          6427 => x"3f7951ff",
          6428 => x"b3933fab",
          6429 => x"3d085482",
          6430 => x"b6980874",
          6431 => x"34805877",
          6432 => x"82b6980c",
          6433 => x"a93d0d04",
          6434 => x"f63d0d7c",
          6435 => x"7e715c71",
          6436 => x"72335759",
          6437 => x"5a5873a0",
          6438 => x"2e098106",
          6439 => x"a2387833",
          6440 => x"78055677",
          6441 => x"76279838",
          6442 => x"8117705b",
          6443 => x"70713356",
          6444 => x"585573a0",
          6445 => x"2e098106",
          6446 => x"86387575",
          6447 => x"26ea3880",
          6448 => x"54738829",
          6449 => x"82b5f405",
          6450 => x"70085255",
          6451 => x"ffb2b63f",
          6452 => x"82b69808",
          6453 => x"53795274",
          6454 => x"0851ffb5",
          6455 => x"b53f82b6",
          6456 => x"980880c5",
          6457 => x"38841533",
          6458 => x"5574812e",
          6459 => x"88387482",
          6460 => x"2e8838b5",
          6461 => x"39fce63f",
          6462 => x"ac39811a",
          6463 => x"5a8c3dfc",
          6464 => x"1153f805",
          6465 => x"51c5c53f",
          6466 => x"82b69808",
          6467 => x"802e9a38",
          6468 => x"ff1b5378",
          6469 => x"527751fd",
          6470 => x"b13f82b6",
          6471 => x"980881ff",
          6472 => x"06557485",
          6473 => x"38745491",
          6474 => x"39811470",
          6475 => x"81ff0651",
          6476 => x"54827427",
          6477 => x"ff8b3880",
          6478 => x"547382b6",
          6479 => x"980c8c3d",
          6480 => x"0d04d33d",
          6481 => x"0db03d08",
          6482 => x"b23d08b4",
          6483 => x"3d08595f",
          6484 => x"5a800baf",
          6485 => x"3d3482b5",
          6486 => x"f03382b5",
          6487 => x"ec08555b",
          6488 => x"7381cb38",
          6489 => x"7382b5e8",
          6490 => x"33555573",
          6491 => x"83388155",
          6492 => x"76802e81",
          6493 => x"bc388170",
          6494 => x"76065556",
          6495 => x"73802e81",
          6496 => x"ad38a851",
          6497 => x"98863f82",
          6498 => x"b6980882",
          6499 => x"b5ec0c82",
          6500 => x"b6980880",
          6501 => x"2e819238",
          6502 => x"93537652",
          6503 => x"82b69808",
          6504 => x"5180ccfa",
          6505 => x"3f82b698",
          6506 => x"08802e8c",
          6507 => x"3882aed0",
          6508 => x"51ffa4af",
          6509 => x"3f80f739",
          6510 => x"82b69808",
          6511 => x"5b82b5ec",
          6512 => x"085380f8",
          6513 => x"52903d70",
          6514 => x"52548187",
          6515 => x"b73f82b6",
          6516 => x"98085682",
          6517 => x"b6980874",
          6518 => x"2e098106",
          6519 => x"80d03882",
          6520 => x"b6980851",
          6521 => x"ffb09e3f",
          6522 => x"82b69808",
          6523 => x"55800b82",
          6524 => x"b6980825",
          6525 => x"a93882b6",
          6526 => x"9808ff05",
          6527 => x"70175555",
          6528 => x"80743480",
          6529 => x"537481ff",
          6530 => x"06527551",
          6531 => x"f8c23f81",
          6532 => x"1b7081ff",
          6533 => x"065c5493",
          6534 => x"7b278338",
          6535 => x"805b74ff",
          6536 => x"2e098106",
          6537 => x"ff973886",
          6538 => x"397582b5",
          6539 => x"e834768c",
          6540 => x"3882b5ec",
          6541 => x"08802e84",
          6542 => x"38f9d63f",
          6543 => x"8f3d5dec",
          6544 => x"c53f82b6",
          6545 => x"9808982b",
          6546 => x"70982c51",
          6547 => x"5978ff2e",
          6548 => x"ee387881",
          6549 => x"ff0682cd",
          6550 => x"c4337098",
          6551 => x"2b70982c",
          6552 => x"82cdc033",
          6553 => x"70982b70",
          6554 => x"972c7198",
          6555 => x"2c057084",
          6556 => x"2982aba4",
          6557 => x"05700815",
          6558 => x"70335151",
          6559 => x"51515959",
          6560 => x"51595d58",
          6561 => x"81567378",
          6562 => x"2e80e938",
          6563 => x"777427b4",
          6564 => x"38748180",
          6565 => x"0a2981ff",
          6566 => x"0a057098",
          6567 => x"2c515580",
          6568 => x"752480ce",
          6569 => x"38765374",
          6570 => x"527751f6",
          6571 => x"853f82b6",
          6572 => x"980881ff",
          6573 => x"06547380",
          6574 => x"2ed73874",
          6575 => x"82cdc034",
          6576 => x"8156b139",
          6577 => x"7481800a",
          6578 => x"2981800a",
          6579 => x"0570982c",
          6580 => x"7081ff06",
          6581 => x"56515573",
          6582 => x"95269738",
          6583 => x"76537452",
          6584 => x"7751f5ce",
          6585 => x"3f82b698",
          6586 => x"0881ff06",
          6587 => x"5473cc38",
          6588 => x"d3398056",
          6589 => x"75802e80",
          6590 => x"ca38811c",
          6591 => x"557482cd",
          6592 => x"c4347498",
          6593 => x"2b70982c",
          6594 => x"82cdc033",
          6595 => x"70982b70",
          6596 => x"982c7010",
          6597 => x"1170822b",
          6598 => x"82aba811",
          6599 => x"335e5151",
          6600 => x"51575851",
          6601 => x"5574772e",
          6602 => x"098106fe",
          6603 => x"923882ab",
          6604 => x"ac14087d",
          6605 => x"0c800b82",
          6606 => x"cdc43480",
          6607 => x"0b82cdc0",
          6608 => x"34923975",
          6609 => x"82cdc434",
          6610 => x"7582cdc0",
          6611 => x"3478af3d",
          6612 => x"34757d0c",
          6613 => x"7e547395",
          6614 => x"26fde138",
          6615 => x"73842982",
          6616 => x"96b00554",
          6617 => x"73080482",
          6618 => x"cdcc3354",
          6619 => x"737e2efd",
          6620 => x"cb3882cd",
          6621 => x"c8335573",
          6622 => x"7527ab38",
          6623 => x"74982b70",
          6624 => x"982c5155",
          6625 => x"7375249e",
          6626 => x"38741a54",
          6627 => x"73338115",
          6628 => x"34748180",
          6629 => x"0a2981ff",
          6630 => x"0a057098",
          6631 => x"2c82cdcc",
          6632 => x"33565155",
          6633 => x"df3982cd",
          6634 => x"cc338111",
          6635 => x"56547482",
          6636 => x"cdcc3473",
          6637 => x"1a54ae3d",
          6638 => x"33743482",
          6639 => x"cdc83354",
          6640 => x"737e2589",
          6641 => x"38811454",
          6642 => x"7382cdc8",
          6643 => x"3482cdcc",
          6644 => x"33708180",
          6645 => x"0a2981ff",
          6646 => x"0a057098",
          6647 => x"2c82cdc8",
          6648 => x"335a5156",
          6649 => x"56747725",
          6650 => x"a83882cd",
          6651 => x"ec085274",
          6652 => x"1a703352",
          6653 => x"54ffa3ba",
          6654 => x"3f748180",
          6655 => x"0a298180",
          6656 => x"0a057098",
          6657 => x"2c82cdc8",
          6658 => x"33565155",
          6659 => x"737524da",
          6660 => x"3882cdcc",
          6661 => x"3370982b",
          6662 => x"70982c82",
          6663 => x"cdc8335a",
          6664 => x"51565674",
          6665 => x"7725fc94",
          6666 => x"3882cdec",
          6667 => x"08528851",
          6668 => x"ffa2ff3f",
          6669 => x"7481800a",
          6670 => x"2981800a",
          6671 => x"0570982c",
          6672 => x"82cdc833",
          6673 => x"56515573",
          6674 => x"7524de38",
          6675 => x"fbee3983",
          6676 => x"7a34800b",
          6677 => x"811b3482",
          6678 => x"cdcc5380",
          6679 => x"52829eec",
          6680 => x"51f39c3f",
          6681 => x"81fd3982",
          6682 => x"cdcc3370",
          6683 => x"81ff0655",
          6684 => x"5573802e",
          6685 => x"fbc63882",
          6686 => x"cdc833ff",
          6687 => x"05547382",
          6688 => x"cdc834ff",
          6689 => x"15547382",
          6690 => x"cdcc3482",
          6691 => x"cdec0852",
          6692 => x"8851ffa2",
          6693 => x"9d3f82cd",
          6694 => x"cc337098",
          6695 => x"2b70982c",
          6696 => x"82cdc833",
          6697 => x"57515657",
          6698 => x"747425ad",
          6699 => x"38741a54",
          6700 => x"81143374",
          6701 => x"3482cdec",
          6702 => x"08527333",
          6703 => x"51ffa1f2",
          6704 => x"3f748180",
          6705 => x"0a298180",
          6706 => x"0a057098",
          6707 => x"2c82cdc8",
          6708 => x"33585155",
          6709 => x"757524d5",
          6710 => x"3882cdec",
          6711 => x"0852a051",
          6712 => x"ffa1cf3f",
          6713 => x"82cdcc33",
          6714 => x"70982b70",
          6715 => x"982c82cd",
          6716 => x"c8335751",
          6717 => x"56577474",
          6718 => x"24fac138",
          6719 => x"82cdec08",
          6720 => x"528851ff",
          6721 => x"a1ac3f74",
          6722 => x"81800a29",
          6723 => x"81800a05",
          6724 => x"70982c82",
          6725 => x"cdc83358",
          6726 => x"51557575",
          6727 => x"25de38fa",
          6728 => x"9b3982cd",
          6729 => x"c8337a05",
          6730 => x"54807434",
          6731 => x"82cdec08",
          6732 => x"528a51ff",
          6733 => x"a0fc3f82",
          6734 => x"cdc85279",
          6735 => x"51f6c93f",
          6736 => x"82b69808",
          6737 => x"81ff0654",
          6738 => x"73963882",
          6739 => x"cdc83354",
          6740 => x"73802e8f",
          6741 => x"38815373",
          6742 => x"527951f1",
          6743 => x"f33f8439",
          6744 => x"807a3480",
          6745 => x"0b82cdcc",
          6746 => x"34800b82",
          6747 => x"cdc83479",
          6748 => x"82b6980c",
          6749 => x"af3d0d04",
          6750 => x"82cdcc33",
          6751 => x"5473802e",
          6752 => x"f9ba3882",
          6753 => x"cdec0852",
          6754 => x"8851ffa0",
          6755 => x"a53f82cd",
          6756 => x"cc33ff05",
          6757 => x"547382cd",
          6758 => x"cc347381",
          6759 => x"ff0654dd",
          6760 => x"3982cdcc",
          6761 => x"3382cdc8",
          6762 => x"33555573",
          6763 => x"752ef98c",
          6764 => x"38ff1454",
          6765 => x"7382cdc8",
          6766 => x"3474982b",
          6767 => x"70982c75",
          6768 => x"81ff0656",
          6769 => x"51557474",
          6770 => x"25ad3874",
          6771 => x"1a548114",
          6772 => x"33743482",
          6773 => x"cdec0852",
          6774 => x"733351ff",
          6775 => x"9fd43f74",
          6776 => x"81800a29",
          6777 => x"81800a05",
          6778 => x"70982c82",
          6779 => x"cdc83358",
          6780 => x"51557575",
          6781 => x"24d53882",
          6782 => x"cdec0852",
          6783 => x"a051ff9f",
          6784 => x"b13f82cd",
          6785 => x"cc337098",
          6786 => x"2b70982c",
          6787 => x"82cdc833",
          6788 => x"57515657",
          6789 => x"747424f8",
          6790 => x"a33882cd",
          6791 => x"ec085288",
          6792 => x"51ff9f8e",
          6793 => x"3f748180",
          6794 => x"0a298180",
          6795 => x"0a057098",
          6796 => x"2c82cdc8",
          6797 => x"33585155",
          6798 => x"757525de",
          6799 => x"38f7fd39",
          6800 => x"82cdcc33",
          6801 => x"7081ff06",
          6802 => x"82cdc833",
          6803 => x"59565474",
          6804 => x"7727f7e8",
          6805 => x"3882cdec",
          6806 => x"08528114",
          6807 => x"547382cd",
          6808 => x"cc34741a",
          6809 => x"70335254",
          6810 => x"ff9ec73f",
          6811 => x"82cdcc33",
          6812 => x"7081ff06",
          6813 => x"82cdc833",
          6814 => x"58565475",
          6815 => x"7526d638",
          6816 => x"f7ba3982",
          6817 => x"cdcc5380",
          6818 => x"52829eec",
          6819 => x"51eef03f",
          6820 => x"800b82cd",
          6821 => x"cc34800b",
          6822 => x"82cdc834",
          6823 => x"f79e397a",
          6824 => x"b03882b5",
          6825 => x"e4085574",
          6826 => x"802ea638",
          6827 => x"7451ffa6",
          6828 => x"d43f82b6",
          6829 => x"980882cd",
          6830 => x"c83482b6",
          6831 => x"980881ff",
          6832 => x"06810553",
          6833 => x"74527951",
          6834 => x"ffa89a3f",
          6835 => x"935b81c0",
          6836 => x"397a8429",
          6837 => x"82b59805",
          6838 => x"fc110856",
          6839 => x"5474802e",
          6840 => x"a7387451",
          6841 => x"ffa69e3f",
          6842 => x"82b69808",
          6843 => x"82cdc834",
          6844 => x"82b69808",
          6845 => x"81ff0681",
          6846 => x"05537452",
          6847 => x"7951ffa7",
          6848 => x"e43fff1b",
          6849 => x"5480fa39",
          6850 => x"73085574",
          6851 => x"802ef6ac",
          6852 => x"387451ff",
          6853 => x"a5ef3f99",
          6854 => x"397a932e",
          6855 => x"098106ae",
          6856 => x"3882b598",
          6857 => x"08557480",
          6858 => x"2ea43874",
          6859 => x"51ffa5d5",
          6860 => x"3f82b698",
          6861 => x"0882cdc8",
          6862 => x"3482b698",
          6863 => x"0881ff06",
          6864 => x"81055374",
          6865 => x"527951ff",
          6866 => x"a79b3f80",
          6867 => x"c3397a84",
          6868 => x"2982b59c",
          6869 => x"05700856",
          6870 => x"5474802e",
          6871 => x"ab387451",
          6872 => x"ffa5a23f",
          6873 => x"82b69808",
          6874 => x"82cdc834",
          6875 => x"82b69808",
          6876 => x"81ff0681",
          6877 => x"05537452",
          6878 => x"7951ffa6",
          6879 => x"e83f811b",
          6880 => x"547381ff",
          6881 => x"065b8939",
          6882 => x"7482cdc8",
          6883 => x"34747a34",
          6884 => x"82cdcc53",
          6885 => x"82cdc833",
          6886 => x"527951ec",
          6887 => x"e23ff59c",
          6888 => x"3982cdcc",
          6889 => x"337081ff",
          6890 => x"0682cdc8",
          6891 => x"33595654",
          6892 => x"747727f5",
          6893 => x"873882cd",
          6894 => x"ec085281",
          6895 => x"14547382",
          6896 => x"cdcc3474",
          6897 => x"1a703352",
          6898 => x"54ff9be6",
          6899 => x"3ff4ed39",
          6900 => x"82cdcc33",
          6901 => x"5473802e",
          6902 => x"f4e23882",
          6903 => x"cdec0852",
          6904 => x"8851ff9b",
          6905 => x"cd3f82cd",
          6906 => x"cc33ff05",
          6907 => x"547382cd",
          6908 => x"cc34f4c8",
          6909 => x"39f93d0d",
          6910 => x"83bff40b",
          6911 => x"82b6900c",
          6912 => x"84800b82",
          6913 => x"b68c23a0",
          6914 => x"80538052",
          6915 => x"83bff451",
          6916 => x"ffaad33f",
          6917 => x"82b69008",
          6918 => x"54805877",
          6919 => x"74348157",
          6920 => x"76811534",
          6921 => x"82b69008",
          6922 => x"54778415",
          6923 => x"34768515",
          6924 => x"3482b690",
          6925 => x"08547786",
          6926 => x"15347687",
          6927 => x"153482b6",
          6928 => x"900882b6",
          6929 => x"8c22ff05",
          6930 => x"fe808007",
          6931 => x"7083ffff",
          6932 => x"0670882a",
          6933 => x"58515556",
          6934 => x"74881734",
          6935 => x"73891734",
          6936 => x"82b68c22",
          6937 => x"70882982",
          6938 => x"b6900805",
          6939 => x"f8115155",
          6940 => x"55778215",
          6941 => x"34768315",
          6942 => x"34893d0d",
          6943 => x"04ff3d0d",
          6944 => x"73528151",
          6945 => x"8472278f",
          6946 => x"38fb1283",
          6947 => x"2a821170",
          6948 => x"83ffff06",
          6949 => x"51515170",
          6950 => x"82b6980c",
          6951 => x"833d0d04",
          6952 => x"f93d0d02",
          6953 => x"a6052202",
          6954 => x"8405aa05",
          6955 => x"22710582",
          6956 => x"b6900871",
          6957 => x"832b7111",
          6958 => x"74832b73",
          6959 => x"11703381",
          6960 => x"12337188",
          6961 => x"2b0702a4",
          6962 => x"05ae0522",
          6963 => x"7181ffff",
          6964 => x"06077088",
          6965 => x"2a535152",
          6966 => x"59545b5b",
          6967 => x"57535455",
          6968 => x"71773470",
          6969 => x"81183482",
          6970 => x"b6900814",
          6971 => x"75882a52",
          6972 => x"54708215",
          6973 => x"34748315",
          6974 => x"3482b690",
          6975 => x"08701770",
          6976 => x"33811233",
          6977 => x"71882b07",
          6978 => x"70832b8f",
          6979 => x"fff80651",
          6980 => x"52565271",
          6981 => x"057383ff",
          6982 => x"ff067088",
          6983 => x"2a545451",
          6984 => x"71821234",
          6985 => x"7281ff06",
          6986 => x"53728312",
          6987 => x"3482b690",
          6988 => x"08165671",
          6989 => x"76347281",
          6990 => x"1734893d",
          6991 => x"0d04fb3d",
          6992 => x"0d82b690",
          6993 => x"08028405",
          6994 => x"9e052270",
          6995 => x"832b7211",
          6996 => x"86113387",
          6997 => x"1233718b",
          6998 => x"2b71832b",
          6999 => x"07585b59",
          7000 => x"52555272",
          7001 => x"05841233",
          7002 => x"85133371",
          7003 => x"882b0770",
          7004 => x"882a5456",
          7005 => x"56527084",
          7006 => x"13347385",
          7007 => x"133482b6",
          7008 => x"90087014",
          7009 => x"84113385",
          7010 => x"1233718b",
          7011 => x"2b71832b",
          7012 => x"07565957",
          7013 => x"52720586",
          7014 => x"12338713",
          7015 => x"3371882b",
          7016 => x"0770882a",
          7017 => x"54565652",
          7018 => x"70861334",
          7019 => x"73871334",
          7020 => x"82b69008",
          7021 => x"13703381",
          7022 => x"12337188",
          7023 => x"2b077081",
          7024 => x"ffff0670",
          7025 => x"882a5351",
          7026 => x"53535371",
          7027 => x"73347081",
          7028 => x"1434873d",
          7029 => x"0d04fa3d",
          7030 => x"0d02a205",
          7031 => x"2282b690",
          7032 => x"0871832b",
          7033 => x"71117033",
          7034 => x"81123371",
          7035 => x"882b0770",
          7036 => x"88291570",
          7037 => x"33811233",
          7038 => x"71982b71",
          7039 => x"902b0753",
          7040 => x"5f535552",
          7041 => x"5a565753",
          7042 => x"54718025",
          7043 => x"80f63872",
          7044 => x"51feab3f",
          7045 => x"82b69008",
          7046 => x"70167033",
          7047 => x"81123371",
          7048 => x"8b2b7183",
          7049 => x"2b077411",
          7050 => x"70338112",
          7051 => x"3371882b",
          7052 => x"0770832b",
          7053 => x"8ffff806",
          7054 => x"51525451",
          7055 => x"535a5853",
          7056 => x"72057488",
          7057 => x"2a545272",
          7058 => x"82133473",
          7059 => x"83133482",
          7060 => x"b6900870",
          7061 => x"16703381",
          7062 => x"1233718b",
          7063 => x"2b71832b",
          7064 => x"07565957",
          7065 => x"55720570",
          7066 => x"33811233",
          7067 => x"71882b07",
          7068 => x"7081ffff",
          7069 => x"0670882a",
          7070 => x"57515258",
          7071 => x"52727434",
          7072 => x"71811534",
          7073 => x"883d0d04",
          7074 => x"fb3d0d82",
          7075 => x"b6900802",
          7076 => x"84059e05",
          7077 => x"2270832b",
          7078 => x"72118211",
          7079 => x"33831233",
          7080 => x"718b2b71",
          7081 => x"832b0759",
          7082 => x"5b595256",
          7083 => x"52730571",
          7084 => x"33811333",
          7085 => x"71882b07",
          7086 => x"028c05a2",
          7087 => x"05227107",
          7088 => x"70882a53",
          7089 => x"51535353",
          7090 => x"71733470",
          7091 => x"81143482",
          7092 => x"b6900870",
          7093 => x"15703381",
          7094 => x"1233718b",
          7095 => x"2b71832b",
          7096 => x"07565957",
          7097 => x"52720582",
          7098 => x"12338313",
          7099 => x"3371882b",
          7100 => x"0770882a",
          7101 => x"54555652",
          7102 => x"70821334",
          7103 => x"72831334",
          7104 => x"82b69008",
          7105 => x"14821133",
          7106 => x"83123371",
          7107 => x"882b0782",
          7108 => x"b6980c52",
          7109 => x"54873d0d",
          7110 => x"04f73d0d",
          7111 => x"7b82b690",
          7112 => x"0831832a",
          7113 => x"7083ffff",
          7114 => x"06705357",
          7115 => x"53fda73f",
          7116 => x"82b69008",
          7117 => x"76832b71",
          7118 => x"11821133",
          7119 => x"83123371",
          7120 => x"8b2b7183",
          7121 => x"2b077511",
          7122 => x"70338112",
          7123 => x"3371982b",
          7124 => x"71902b07",
          7125 => x"53424051",
          7126 => x"535b5855",
          7127 => x"59547280",
          7128 => x"258d3882",
          7129 => x"80805275",
          7130 => x"51fe9d3f",
          7131 => x"81843984",
          7132 => x"14338515",
          7133 => x"33718b2b",
          7134 => x"71832b07",
          7135 => x"76117988",
          7136 => x"2a535155",
          7137 => x"58557686",
          7138 => x"14347581",
          7139 => x"ff065675",
          7140 => x"87143482",
          7141 => x"b6900870",
          7142 => x"19841233",
          7143 => x"85133371",
          7144 => x"882b0770",
          7145 => x"882a5457",
          7146 => x"5b565372",
          7147 => x"84163473",
          7148 => x"85163482",
          7149 => x"b6900818",
          7150 => x"53800b86",
          7151 => x"1434800b",
          7152 => x"87143482",
          7153 => x"b6900853",
          7154 => x"76841434",
          7155 => x"75851434",
          7156 => x"82b69008",
          7157 => x"18703381",
          7158 => x"12337188",
          7159 => x"2b077082",
          7160 => x"80800770",
          7161 => x"882a5351",
          7162 => x"55565474",
          7163 => x"74347281",
          7164 => x"15348b3d",
          7165 => x"0d04ff3d",
          7166 => x"0d735282",
          7167 => x"b6900884",
          7168 => x"38f7f23f",
          7169 => x"71802e86",
          7170 => x"387151fe",
          7171 => x"8c3f833d",
          7172 => x"0d04f53d",
          7173 => x"0d807e52",
          7174 => x"58f8e23f",
          7175 => x"82b69808",
          7176 => x"83ffff06",
          7177 => x"82b69008",
          7178 => x"84113385",
          7179 => x"12337188",
          7180 => x"2b07705f",
          7181 => x"5956585a",
          7182 => x"81ffff59",
          7183 => x"75782e80",
          7184 => x"cb387588",
          7185 => x"29177033",
          7186 => x"81123371",
          7187 => x"882b0770",
          7188 => x"81ffff06",
          7189 => x"79317083",
          7190 => x"ffff0670",
          7191 => x"7f275253",
          7192 => x"51565955",
          7193 => x"7779278a",
          7194 => x"3873802e",
          7195 => x"85387578",
          7196 => x"5a5b8415",
          7197 => x"33851633",
          7198 => x"71882b07",
          7199 => x"575475c2",
          7200 => x"387881ff",
          7201 => x"ff2e8538",
          7202 => x"7a795956",
          7203 => x"8076832b",
          7204 => x"82b69008",
          7205 => x"11703381",
          7206 => x"12337188",
          7207 => x"2b077081",
          7208 => x"ffff0651",
          7209 => x"525a565c",
          7210 => x"5573752e",
          7211 => x"83388155",
          7212 => x"80547978",
          7213 => x"2681cc38",
          7214 => x"74547480",
          7215 => x"2e81c438",
          7216 => x"777a2e09",
          7217 => x"81068938",
          7218 => x"7551f8f2",
          7219 => x"3f81ac39",
          7220 => x"82808053",
          7221 => x"79527551",
          7222 => x"f7c63f82",
          7223 => x"b6900870",
          7224 => x"1c861133",
          7225 => x"87123371",
          7226 => x"8b2b7183",
          7227 => x"2b07535a",
          7228 => x"5e557405",
          7229 => x"7a177083",
          7230 => x"ffff0670",
          7231 => x"882a5c59",
          7232 => x"56547884",
          7233 => x"15347681",
          7234 => x"ff065776",
          7235 => x"85153482",
          7236 => x"b6900875",
          7237 => x"832b7111",
          7238 => x"721e8611",
          7239 => x"33871233",
          7240 => x"71882b07",
          7241 => x"70882a53",
          7242 => x"5b5e535a",
          7243 => x"56547386",
          7244 => x"19347587",
          7245 => x"193482b6",
          7246 => x"9008701c",
          7247 => x"84113385",
          7248 => x"1233718b",
          7249 => x"2b71832b",
          7250 => x"07535d5a",
          7251 => x"55740554",
          7252 => x"78861534",
          7253 => x"76871534",
          7254 => x"82b69008",
          7255 => x"7016711d",
          7256 => x"84113385",
          7257 => x"12337188",
          7258 => x"2b077088",
          7259 => x"2a535a5f",
          7260 => x"52565473",
          7261 => x"84163475",
          7262 => x"85163482",
          7263 => x"b690081b",
          7264 => x"84055473",
          7265 => x"82b6980c",
          7266 => x"8d3d0d04",
          7267 => x"fe3d0d74",
          7268 => x"5282b690",
          7269 => x"088438f4",
          7270 => x"dc3f7153",
          7271 => x"71802e8b",
          7272 => x"387151fc",
          7273 => x"ed3f82b6",
          7274 => x"98085372",
          7275 => x"82b6980c",
          7276 => x"843d0d04",
          7277 => x"ee3d0d64",
          7278 => x"66405c80",
          7279 => x"70424082",
          7280 => x"b6900860",
          7281 => x"2e098106",
          7282 => x"8438f4a9",
          7283 => x"3f7b8e38",
          7284 => x"7e51ffb8",
          7285 => x"3f82b698",
          7286 => x"085483c7",
          7287 => x"397e8b38",
          7288 => x"7b51fc92",
          7289 => x"3f7e5483",
          7290 => x"ba397e51",
          7291 => x"f58f3f82",
          7292 => x"b6980883",
          7293 => x"ffff0682",
          7294 => x"b690087d",
          7295 => x"7131832a",
          7296 => x"7083ffff",
          7297 => x"0670832b",
          7298 => x"73117033",
          7299 => x"81123371",
          7300 => x"882b0770",
          7301 => x"75317083",
          7302 => x"ffff0670",
          7303 => x"8829fc05",
          7304 => x"7388291a",
          7305 => x"70338112",
          7306 => x"3371882b",
          7307 => x"0770902b",
          7308 => x"53444e53",
          7309 => x"4841525c",
          7310 => x"545b415c",
          7311 => x"565b5b73",
          7312 => x"80258f38",
          7313 => x"7681ffff",
          7314 => x"06753170",
          7315 => x"83ffff06",
          7316 => x"42548216",
          7317 => x"33831733",
          7318 => x"71882b07",
          7319 => x"7088291c",
          7320 => x"70338112",
          7321 => x"3371982b",
          7322 => x"71902b07",
          7323 => x"53474552",
          7324 => x"56547380",
          7325 => x"258b3878",
          7326 => x"75317083",
          7327 => x"ffff0641",
          7328 => x"54777b27",
          7329 => x"81fe3860",
          7330 => x"1854737b",
          7331 => x"2e098106",
          7332 => x"8f387851",
          7333 => x"f6c03f7a",
          7334 => x"83ffff06",
          7335 => x"5881e539",
          7336 => x"7f8e387a",
          7337 => x"74248938",
          7338 => x"7851f6aa",
          7339 => x"3f81a539",
          7340 => x"7f18557a",
          7341 => x"752480c8",
          7342 => x"38791d82",
          7343 => x"11338312",
          7344 => x"3371882b",
          7345 => x"07535754",
          7346 => x"f4f43f80",
          7347 => x"527851f7",
          7348 => x"b73f82b6",
          7349 => x"980883ff",
          7350 => x"ff067e54",
          7351 => x"7c537083",
          7352 => x"2b82b690",
          7353 => x"08118405",
          7354 => x"535559ff",
          7355 => x"93ad3f82",
          7356 => x"b6900814",
          7357 => x"84057583",
          7358 => x"ffff0659",
          7359 => x"5c818539",
          7360 => x"6015547a",
          7361 => x"742480d4",
          7362 => x"387851f5",
          7363 => x"c93f82b6",
          7364 => x"90081d82",
          7365 => x"11338312",
          7366 => x"3371882b",
          7367 => x"07534354",
          7368 => x"f49c3f80",
          7369 => x"527851f6",
          7370 => x"df3f82b6",
          7371 => x"980883ff",
          7372 => x"ff067e54",
          7373 => x"7c537083",
          7374 => x"2b82b690",
          7375 => x"08118405",
          7376 => x"535559ff",
          7377 => x"92d53f82",
          7378 => x"b6900814",
          7379 => x"84056062",
          7380 => x"0519555c",
          7381 => x"7383ffff",
          7382 => x"0658a939",
          7383 => x"7b7f5254",
          7384 => x"f9b03f82",
          7385 => x"b698085c",
          7386 => x"82b69808",
          7387 => x"802e9338",
          7388 => x"7d537352",
          7389 => x"82b69808",
          7390 => x"51ff96e9",
          7391 => x"3f7351f7",
          7392 => x"983f7a58",
          7393 => x"7a782799",
          7394 => x"3880537a",
          7395 => x"527851f2",
          7396 => x"8f3f7a19",
          7397 => x"832b82b6",
          7398 => x"90080584",
          7399 => x"0551f6f9",
          7400 => x"3f7b5473",
          7401 => x"82b6980c",
          7402 => x"943d0d04",
          7403 => x"fc3d0d77",
          7404 => x"77297052",
          7405 => x"54fbd53f",
          7406 => x"82b69808",
          7407 => x"5582b698",
          7408 => x"08802e8e",
          7409 => x"38735380",
          7410 => x"5282b698",
          7411 => x"0851ff9b",
          7412 => x"953f7482",
          7413 => x"b6980c86",
          7414 => x"3d0d04ff",
          7415 => x"3d0d028f",
          7416 => x"05335181",
          7417 => x"52707226",
          7418 => x"873882b6",
          7419 => x"94113352",
          7420 => x"7182b698",
          7421 => x"0c833d0d",
          7422 => x"04fc3d0d",
          7423 => x"029b0533",
          7424 => x"0284059f",
          7425 => x"05335653",
          7426 => x"83517281",
          7427 => x"2680e038",
          7428 => x"72842b87",
          7429 => x"c0928c11",
          7430 => x"53518854",
          7431 => x"74802e84",
          7432 => x"38818854",
          7433 => x"73720c87",
          7434 => x"c0928c11",
          7435 => x"5181710c",
          7436 => x"850b87c0",
          7437 => x"988c0c70",
          7438 => x"52710870",
          7439 => x"82065151",
          7440 => x"70802e8a",
          7441 => x"3887c098",
          7442 => x"8c085170",
          7443 => x"ec387108",
          7444 => x"fc808006",
          7445 => x"52719238",
          7446 => x"87c0988c",
          7447 => x"08517080",
          7448 => x"2e873871",
          7449 => x"82b69414",
          7450 => x"3482b694",
          7451 => x"13335170",
          7452 => x"82b6980c",
          7453 => x"863d0d04",
          7454 => x"f33d0d60",
          7455 => x"6264028c",
          7456 => x"05bf0533",
          7457 => x"5740585b",
          7458 => x"8374525a",
          7459 => x"fecd3f82",
          7460 => x"b6980881",
          7461 => x"067a5452",
          7462 => x"7181be38",
          7463 => x"71727584",
          7464 => x"2b87c092",
          7465 => x"801187c0",
          7466 => x"928c1287",
          7467 => x"c0928413",
          7468 => x"415a4057",
          7469 => x"5a58850b",
          7470 => x"87c0988c",
          7471 => x"0c767d0c",
          7472 => x"84760c75",
          7473 => x"0870852a",
          7474 => x"70810651",
          7475 => x"53547180",
          7476 => x"2e8e387b",
          7477 => x"0852717b",
          7478 => x"7081055d",
          7479 => x"34811959",
          7480 => x"8074a206",
          7481 => x"53537173",
          7482 => x"2e833881",
          7483 => x"537883ff",
          7484 => x"268f3872",
          7485 => x"802e8a38",
          7486 => x"87c0988c",
          7487 => x"085271c3",
          7488 => x"3887c098",
          7489 => x"8c085271",
          7490 => x"802e8738",
          7491 => x"7884802e",
          7492 => x"99388176",
          7493 => x"0c87c092",
          7494 => x"8c155372",
          7495 => x"08708206",
          7496 => x"515271f7",
          7497 => x"38ff1a5a",
          7498 => x"8d398480",
          7499 => x"17811970",
          7500 => x"81ff065a",
          7501 => x"53577980",
          7502 => x"2e903873",
          7503 => x"fc808006",
          7504 => x"52718738",
          7505 => x"7d7826fe",
          7506 => x"ed3873fc",
          7507 => x"80800652",
          7508 => x"71802e83",
          7509 => x"38815271",
          7510 => x"537282b6",
          7511 => x"980c8f3d",
          7512 => x"0d04f33d",
          7513 => x"0d606264",
          7514 => x"028c05bf",
          7515 => x"05335740",
          7516 => x"585b8359",
          7517 => x"80745258",
          7518 => x"fce13f82",
          7519 => x"b6980881",
          7520 => x"06795452",
          7521 => x"71782e09",
          7522 => x"810681b1",
          7523 => x"38777484",
          7524 => x"2b87c092",
          7525 => x"801187c0",
          7526 => x"928c1287",
          7527 => x"c0928413",
          7528 => x"40595f56",
          7529 => x"5a850b87",
          7530 => x"c0988c0c",
          7531 => x"767d0c82",
          7532 => x"760c8058",
          7533 => x"75087084",
          7534 => x"2a708106",
          7535 => x"51535471",
          7536 => x"802e8c38",
          7537 => x"7a708105",
          7538 => x"5c337c0c",
          7539 => x"81185873",
          7540 => x"812a7081",
          7541 => x"06515271",
          7542 => x"802e8a38",
          7543 => x"87c0988c",
          7544 => x"085271d0",
          7545 => x"3887c098",
          7546 => x"8c085271",
          7547 => x"802e8738",
          7548 => x"7784802e",
          7549 => x"99388176",
          7550 => x"0c87c092",
          7551 => x"8c155372",
          7552 => x"08708206",
          7553 => x"515271f7",
          7554 => x"38ff1959",
          7555 => x"8d39811a",
          7556 => x"7081ff06",
          7557 => x"84801959",
          7558 => x"5b527880",
          7559 => x"2e903873",
          7560 => x"fc808006",
          7561 => x"52718738",
          7562 => x"7d7a26fe",
          7563 => x"f83873fc",
          7564 => x"80800652",
          7565 => x"71802e83",
          7566 => x"38815271",
          7567 => x"537282b6",
          7568 => x"980c8f3d",
          7569 => x"0d04fa3d",
          7570 => x"0d7a0284",
          7571 => x"05a30533",
          7572 => x"028805a7",
          7573 => x"05337154",
          7574 => x"545657fa",
          7575 => x"fe3f82b6",
          7576 => x"98088106",
          7577 => x"53835472",
          7578 => x"80fe3885",
          7579 => x"0b87c098",
          7580 => x"8c0c8156",
          7581 => x"71762e80",
          7582 => x"dc387176",
          7583 => x"24933874",
          7584 => x"842b87c0",
          7585 => x"928c1154",
          7586 => x"5471802e",
          7587 => x"8d3880d4",
          7588 => x"3971832e",
          7589 => x"80c63880",
          7590 => x"cb397208",
          7591 => x"70812a70",
          7592 => x"81065151",
          7593 => x"5271802e",
          7594 => x"8a3887c0",
          7595 => x"988c0852",
          7596 => x"71e83887",
          7597 => x"c0988c08",
          7598 => x"52719638",
          7599 => x"81730c87",
          7600 => x"c0928c14",
          7601 => x"53720870",
          7602 => x"82065152",
          7603 => x"71f73896",
          7604 => x"39805692",
          7605 => x"3988800a",
          7606 => x"770c8539",
          7607 => x"8180770c",
          7608 => x"72568339",
          7609 => x"84567554",
          7610 => x"7382b698",
          7611 => x"0c883d0d",
          7612 => x"04fe3d0d",
          7613 => x"74811133",
          7614 => x"71337188",
          7615 => x"2b0782b6",
          7616 => x"980c5351",
          7617 => x"843d0d04",
          7618 => x"fd3d0d75",
          7619 => x"83113382",
          7620 => x"12337190",
          7621 => x"2b71882b",
          7622 => x"07811433",
          7623 => x"70720788",
          7624 => x"2b753371",
          7625 => x"0782b698",
          7626 => x"0c525354",
          7627 => x"56545285",
          7628 => x"3d0d04ff",
          7629 => x"3d0d7302",
          7630 => x"84059205",
          7631 => x"22525270",
          7632 => x"72708105",
          7633 => x"54347088",
          7634 => x"2a517072",
          7635 => x"34833d0d",
          7636 => x"04ff3d0d",
          7637 => x"73755252",
          7638 => x"70727081",
          7639 => x"05543470",
          7640 => x"882a5170",
          7641 => x"72708105",
          7642 => x"54347088",
          7643 => x"2a517072",
          7644 => x"70810554",
          7645 => x"3470882a",
          7646 => x"51707234",
          7647 => x"833d0d04",
          7648 => x"fe3d0d76",
          7649 => x"75775454",
          7650 => x"5170802e",
          7651 => x"92387170",
          7652 => x"81055333",
          7653 => x"73708105",
          7654 => x"5534ff11",
          7655 => x"51eb3984",
          7656 => x"3d0d04fe",
          7657 => x"3d0d7577",
          7658 => x"76545253",
          7659 => x"72727081",
          7660 => x"055434ff",
          7661 => x"115170f4",
          7662 => x"38843d0d",
          7663 => x"04fc3d0d",
          7664 => x"78777956",
          7665 => x"56537470",
          7666 => x"81055633",
          7667 => x"74708105",
          7668 => x"56337171",
          7669 => x"31ff1656",
          7670 => x"52525272",
          7671 => x"802e8638",
          7672 => x"71802ee2",
          7673 => x"387182b6",
          7674 => x"980c863d",
          7675 => x"0d04fe3d",
          7676 => x"0d747654",
          7677 => x"51893971",
          7678 => x"732e8a38",
          7679 => x"81115170",
          7680 => x"335271f3",
          7681 => x"38703382",
          7682 => x"b6980c84",
          7683 => x"3d0d0480",
          7684 => x"0b82b698",
          7685 => x"0c04800b",
          7686 => x"82b6980c",
          7687 => x"04f73d0d",
          7688 => x"7b56800b",
          7689 => x"83173356",
          7690 => x"5a747a2e",
          7691 => x"80d63881",
          7692 => x"54b01608",
          7693 => x"53b41670",
          7694 => x"53811733",
          7695 => x"5259faa2",
          7696 => x"3f82b698",
          7697 => x"087a2e09",
          7698 => x"8106b738",
          7699 => x"82b69808",
          7700 => x"831734b0",
          7701 => x"160870a4",
          7702 => x"1808319c",
          7703 => x"18085956",
          7704 => x"58747727",
          7705 => x"9f388216",
          7706 => x"33557482",
          7707 => x"2e098106",
          7708 => x"93388154",
          7709 => x"76185378",
          7710 => x"52811633",
          7711 => x"51f9e33f",
          7712 => x"8339815a",
          7713 => x"7982b698",
          7714 => x"0c8b3d0d",
          7715 => x"04fa3d0d",
          7716 => x"787a5656",
          7717 => x"805774b0",
          7718 => x"17082eaf",
          7719 => x"387551fe",
          7720 => x"fc3f82b6",
          7721 => x"98085782",
          7722 => x"b698089f",
          7723 => x"38815474",
          7724 => x"53b41652",
          7725 => x"81163351",
          7726 => x"f7be3f82",
          7727 => x"b6980880",
          7728 => x"2e8538ff",
          7729 => x"55815774",
          7730 => x"b0170c76",
          7731 => x"82b6980c",
          7732 => x"883d0d04",
          7733 => x"f83d0d7a",
          7734 => x"705257fe",
          7735 => x"c03f82b6",
          7736 => x"98085882",
          7737 => x"b6980881",
          7738 => x"91387633",
          7739 => x"5574832e",
          7740 => x"09810680",
          7741 => x"f0388417",
          7742 => x"33597881",
          7743 => x"2e098106",
          7744 => x"80e33884",
          7745 => x"805382b6",
          7746 => x"980852b4",
          7747 => x"17705256",
          7748 => x"fd913f82",
          7749 => x"d4d55284",
          7750 => x"b21751fc",
          7751 => x"963f848b",
          7752 => x"85a4d252",
          7753 => x"7551fca9",
          7754 => x"3f868a85",
          7755 => x"e4f25284",
          7756 => x"981751fc",
          7757 => x"9c3f9017",
          7758 => x"0852849c",
          7759 => x"1751fc91",
          7760 => x"3f8c1708",
          7761 => x"5284a017",
          7762 => x"51fc863f",
          7763 => x"a0170881",
          7764 => x"0570b019",
          7765 => x"0c795553",
          7766 => x"75528117",
          7767 => x"3351f882",
          7768 => x"3f778418",
          7769 => x"34805380",
          7770 => x"52811733",
          7771 => x"51f9d73f",
          7772 => x"82b69808",
          7773 => x"802e8338",
          7774 => x"81587782",
          7775 => x"b6980c8a",
          7776 => x"3d0d04fb",
          7777 => x"3d0d77fe",
          7778 => x"1a981208",
          7779 => x"fe055556",
          7780 => x"54805674",
          7781 => x"73278d38",
          7782 => x"8a142275",
          7783 => x"7129ac16",
          7784 => x"08055753",
          7785 => x"7582b698",
          7786 => x"0c873d0d",
          7787 => x"04f93d0d",
          7788 => x"7a7a7008",
          7789 => x"56545781",
          7790 => x"772781df",
          7791 => x"38769815",
          7792 => x"082781d7",
          7793 => x"38ff7433",
          7794 => x"54587282",
          7795 => x"2e80f538",
          7796 => x"72822489",
          7797 => x"3872812e",
          7798 => x"8d3881bf",
          7799 => x"3972832e",
          7800 => x"818e3881",
          7801 => x"b6397681",
          7802 => x"2a177089",
          7803 => x"2aa41608",
          7804 => x"05537452",
          7805 => x"55fd963f",
          7806 => x"82b69808",
          7807 => x"819f3874",
          7808 => x"83ff0614",
          7809 => x"b4113381",
          7810 => x"1770892a",
          7811 => x"a4180805",
          7812 => x"55765457",
          7813 => x"5753fcf5",
          7814 => x"3f82b698",
          7815 => x"0880fe38",
          7816 => x"7483ff06",
          7817 => x"14b41133",
          7818 => x"70882b78",
          7819 => x"07798106",
          7820 => x"71842a5c",
          7821 => x"52585153",
          7822 => x"7280e238",
          7823 => x"759fff06",
          7824 => x"5880da39",
          7825 => x"76882aa4",
          7826 => x"15080552",
          7827 => x"7351fcbd",
          7828 => x"3f82b698",
          7829 => x"0880c638",
          7830 => x"761083fe",
          7831 => x"067405b4",
          7832 => x"0551f98d",
          7833 => x"3f82b698",
          7834 => x"0883ffff",
          7835 => x"0658ae39",
          7836 => x"76872aa4",
          7837 => x"15080552",
          7838 => x"7351fc91",
          7839 => x"3f82b698",
          7840 => x"089b3876",
          7841 => x"822b83fc",
          7842 => x"067405b4",
          7843 => x"0551f8f8",
          7844 => x"3f82b698",
          7845 => x"08f00a06",
          7846 => x"58833981",
          7847 => x"587782b6",
          7848 => x"980c893d",
          7849 => x"0d04f83d",
          7850 => x"0d7a7c7e",
          7851 => x"5a585682",
          7852 => x"59817727",
          7853 => x"829e3876",
          7854 => x"98170827",
          7855 => x"82963875",
          7856 => x"33537279",
          7857 => x"2e819d38",
          7858 => x"72792489",
          7859 => x"3872812e",
          7860 => x"8d388280",
          7861 => x"3972832e",
          7862 => x"81b83881",
          7863 => x"f7397681",
          7864 => x"2a177089",
          7865 => x"2aa41808",
          7866 => x"05537652",
          7867 => x"55fb9e3f",
          7868 => x"82b69808",
          7869 => x"5982b698",
          7870 => x"0881d938",
          7871 => x"7483ff06",
          7872 => x"16b40581",
          7873 => x"16788106",
          7874 => x"59565477",
          7875 => x"5376802e",
          7876 => x"8f387784",
          7877 => x"2b9ff006",
          7878 => x"74338f06",
          7879 => x"71075153",
          7880 => x"72743481",
          7881 => x"0b831734",
          7882 => x"74892aa4",
          7883 => x"17080552",
          7884 => x"7551fad9",
          7885 => x"3f82b698",
          7886 => x"085982b6",
          7887 => x"98088194",
          7888 => x"387483ff",
          7889 => x"0616b405",
          7890 => x"78842a54",
          7891 => x"54768f38",
          7892 => x"77882a74",
          7893 => x"3381f006",
          7894 => x"718f0607",
          7895 => x"51537274",
          7896 => x"3480ec39",
          7897 => x"76882aa4",
          7898 => x"17080552",
          7899 => x"7551fa9d",
          7900 => x"3f82b698",
          7901 => x"085982b6",
          7902 => x"980880d8",
          7903 => x"387783ff",
          7904 => x"ff065276",
          7905 => x"1083fe06",
          7906 => x"7605b405",
          7907 => x"51f7a43f",
          7908 => x"be397687",
          7909 => x"2aa41708",
          7910 => x"05527551",
          7911 => x"f9ef3f82",
          7912 => x"b6980859",
          7913 => x"82b69808",
          7914 => x"ab3877f0",
          7915 => x"0a067782",
          7916 => x"2b83fc06",
          7917 => x"7018b405",
          7918 => x"70545154",
          7919 => x"54f6c93f",
          7920 => x"82b69808",
          7921 => x"8f0a0674",
          7922 => x"07527251",
          7923 => x"f7833f81",
          7924 => x"0b831734",
          7925 => x"7882b698",
          7926 => x"0c8a3d0d",
          7927 => x"04f83d0d",
          7928 => x"7a7c7e72",
          7929 => x"08595656",
          7930 => x"59817527",
          7931 => x"a4387498",
          7932 => x"1708279d",
          7933 => x"3873802e",
          7934 => x"aa38ff53",
          7935 => x"73527551",
          7936 => x"fda43f82",
          7937 => x"b6980854",
          7938 => x"82b69808",
          7939 => x"80f23893",
          7940 => x"39825480",
          7941 => x"eb398154",
          7942 => x"80e63982",
          7943 => x"b6980854",
          7944 => x"80de3974",
          7945 => x"527851fb",
          7946 => x"843f82b6",
          7947 => x"98085882",
          7948 => x"b6980880",
          7949 => x"2e80c738",
          7950 => x"82b69808",
          7951 => x"812ed238",
          7952 => x"82b69808",
          7953 => x"ff2ecf38",
          7954 => x"80537452",
          7955 => x"7551fcd6",
          7956 => x"3f82b698",
          7957 => x"08c53898",
          7958 => x"1608fe11",
          7959 => x"90180857",
          7960 => x"55577474",
          7961 => x"27903881",
          7962 => x"1590170c",
          7963 => x"84163381",
          7964 => x"07547384",
          7965 => x"17347755",
          7966 => x"767826ff",
          7967 => x"a6388054",
          7968 => x"7382b698",
          7969 => x"0c8a3d0d",
          7970 => x"04f63d0d",
          7971 => x"7c7e7108",
          7972 => x"595b5b79",
          7973 => x"95388c17",
          7974 => x"08587780",
          7975 => x"2e883898",
          7976 => x"17087826",
          7977 => x"b2388158",
          7978 => x"ae397952",
          7979 => x"7a51f9fd",
          7980 => x"3f815574",
          7981 => x"82b69808",
          7982 => x"2782e038",
          7983 => x"82b69808",
          7984 => x"5582b698",
          7985 => x"08ff2e82",
          7986 => x"d2389817",
          7987 => x"0882b698",
          7988 => x"082682c7",
          7989 => x"38795890",
          7990 => x"17087056",
          7991 => x"5473802e",
          7992 => x"82b93877",
          7993 => x"7a2e0981",
          7994 => x"0680e238",
          7995 => x"811a5698",
          7996 => x"17087626",
          7997 => x"83388256",
          7998 => x"75527a51",
          7999 => x"f9af3f80",
          8000 => x"5982b698",
          8001 => x"08812e09",
          8002 => x"81068638",
          8003 => x"82b69808",
          8004 => x"5982b698",
          8005 => x"08097030",
          8006 => x"70720780",
          8007 => x"25707c07",
          8008 => x"82b69808",
          8009 => x"54515155",
          8010 => x"557381ef",
          8011 => x"3882b698",
          8012 => x"08802e95",
          8013 => x"388c1708",
          8014 => x"54817427",
          8015 => x"90387398",
          8016 => x"18082789",
          8017 => x"38735885",
          8018 => x"397580db",
          8019 => x"38775681",
          8020 => x"16569817",
          8021 => x"08762689",
          8022 => x"38825675",
          8023 => x"782681ac",
          8024 => x"3875527a",
          8025 => x"51f8c63f",
          8026 => x"82b69808",
          8027 => x"802eb838",
          8028 => x"805982b6",
          8029 => x"9808812e",
          8030 => x"09810686",
          8031 => x"3882b698",
          8032 => x"085982b6",
          8033 => x"98080970",
          8034 => x"30707207",
          8035 => x"8025707c",
          8036 => x"07515155",
          8037 => x"557380f8",
          8038 => x"3875782e",
          8039 => x"098106ff",
          8040 => x"ae387355",
          8041 => x"80f539ff",
          8042 => x"53755276",
          8043 => x"51f9f73f",
          8044 => x"82b69808",
          8045 => x"82b69808",
          8046 => x"307082b6",
          8047 => x"98080780",
          8048 => x"25515555",
          8049 => x"79802e94",
          8050 => x"3873802e",
          8051 => x"8f387553",
          8052 => x"79527651",
          8053 => x"f9d03f82",
          8054 => x"b6980855",
          8055 => x"74a53875",
          8056 => x"8c180c98",
          8057 => x"1708fe05",
          8058 => x"90180856",
          8059 => x"54747426",
          8060 => x"8638ff15",
          8061 => x"90180c84",
          8062 => x"17338107",
          8063 => x"54738418",
          8064 => x"349739ff",
          8065 => x"5674812e",
          8066 => x"90388c39",
          8067 => x"80558c39",
          8068 => x"82b69808",
          8069 => x"55853981",
          8070 => x"56755574",
          8071 => x"82b6980c",
          8072 => x"8c3d0d04",
          8073 => x"f83d0d7a",
          8074 => x"705255f3",
          8075 => x"f03f82b6",
          8076 => x"98085881",
          8077 => x"5682b698",
          8078 => x"0880d838",
          8079 => x"7b527451",
          8080 => x"f6c13f82",
          8081 => x"b6980882",
          8082 => x"b69808b0",
          8083 => x"170c5984",
          8084 => x"80537752",
          8085 => x"b4157052",
          8086 => x"57f2c83f",
          8087 => x"77568439",
          8088 => x"8116568a",
          8089 => x"15225875",
          8090 => x"78279738",
          8091 => x"81547519",
          8092 => x"53765281",
          8093 => x"153351ed",
          8094 => x"e93f82b6",
          8095 => x"9808802e",
          8096 => x"df388a15",
          8097 => x"22763270",
          8098 => x"30707207",
          8099 => x"709f2a53",
          8100 => x"51565675",
          8101 => x"82b6980c",
          8102 => x"8a3d0d04",
          8103 => x"f83d0d7a",
          8104 => x"7c710858",
          8105 => x"565774f0",
          8106 => x"800a2680",
          8107 => x"f138749f",
          8108 => x"06537280",
          8109 => x"e9387490",
          8110 => x"180c8817",
          8111 => x"085473aa",
          8112 => x"38753353",
          8113 => x"82732788",
          8114 => x"38a81608",
          8115 => x"54739b38",
          8116 => x"74852a53",
          8117 => x"820b8817",
          8118 => x"225a5872",
          8119 => x"792780fe",
          8120 => x"38a81608",
          8121 => x"98180c80",
          8122 => x"cd398a16",
          8123 => x"2270892b",
          8124 => x"54587275",
          8125 => x"26b23873",
          8126 => x"527651f5",
          8127 => x"b03f82b6",
          8128 => x"98085482",
          8129 => x"b69808ff",
          8130 => x"2ebd3881",
          8131 => x"0b82b698",
          8132 => x"08278b38",
          8133 => x"98160882",
          8134 => x"b6980826",
          8135 => x"85388258",
          8136 => x"bd397473",
          8137 => x"3155cb39",
          8138 => x"73527551",
          8139 => x"f4d53f82",
          8140 => x"b6980898",
          8141 => x"180c7394",
          8142 => x"180c9817",
          8143 => x"08538258",
          8144 => x"72802e9a",
          8145 => x"38853981",
          8146 => x"58943974",
          8147 => x"892a1398",
          8148 => x"180c7483",
          8149 => x"ff0616b4",
          8150 => x"059c180c",
          8151 => x"80587782",
          8152 => x"b6980c8a",
          8153 => x"3d0d04f8",
          8154 => x"3d0d7a70",
          8155 => x"08901208",
          8156 => x"a0055957",
          8157 => x"54f0800a",
          8158 => x"77278638",
          8159 => x"800b9815",
          8160 => x"0c981408",
          8161 => x"53845572",
          8162 => x"802e81cb",
          8163 => x"387683ff",
          8164 => x"06587781",
          8165 => x"b5388113",
          8166 => x"98150c94",
          8167 => x"14085574",
          8168 => x"92387685",
          8169 => x"2a881722",
          8170 => x"56537473",
          8171 => x"26819b38",
          8172 => x"80c0398a",
          8173 => x"1622ff05",
          8174 => x"77892a06",
          8175 => x"5372818a",
          8176 => x"38745273",
          8177 => x"51f3e63f",
          8178 => x"82b69808",
          8179 => x"53825581",
          8180 => x"0b82b698",
          8181 => x"082780ff",
          8182 => x"38815582",
          8183 => x"b69808ff",
          8184 => x"2e80f438",
          8185 => x"98160882",
          8186 => x"b6980826",
          8187 => x"80ca387b",
          8188 => x"8a387798",
          8189 => x"150c8455",
          8190 => x"80dd3994",
          8191 => x"14085273",
          8192 => x"51f9863f",
          8193 => x"82b69808",
          8194 => x"53875582",
          8195 => x"b6980880",
          8196 => x"2e80c438",
          8197 => x"825582b6",
          8198 => x"9808812e",
          8199 => x"ba388155",
          8200 => x"82b69808",
          8201 => x"ff2eb038",
          8202 => x"82b69808",
          8203 => x"527551fb",
          8204 => x"f33f82b6",
          8205 => x"9808a038",
          8206 => x"7294150c",
          8207 => x"72527551",
          8208 => x"f2c13f82",
          8209 => x"b6980898",
          8210 => x"150c7690",
          8211 => x"150c7716",
          8212 => x"b4059c15",
          8213 => x"0c805574",
          8214 => x"82b6980c",
          8215 => x"8a3d0d04",
          8216 => x"f73d0d7b",
          8217 => x"7d71085b",
          8218 => x"5b578052",
          8219 => x"7651fcac",
          8220 => x"3f82b698",
          8221 => x"085482b6",
          8222 => x"980880ec",
          8223 => x"3882b698",
          8224 => x"08569817",
          8225 => x"08527851",
          8226 => x"f0833f82",
          8227 => x"b6980854",
          8228 => x"82b69808",
          8229 => x"80d23882",
          8230 => x"b698089c",
          8231 => x"18087033",
          8232 => x"51545872",
          8233 => x"81e52e09",
          8234 => x"81068338",
          8235 => x"815882b6",
          8236 => x"98085572",
          8237 => x"83388155",
          8238 => x"77750753",
          8239 => x"72802e8e",
          8240 => x"38811656",
          8241 => x"757a2e09",
          8242 => x"81068838",
          8243 => x"a53982b6",
          8244 => x"98085681",
          8245 => x"527651fd",
          8246 => x"8e3f82b6",
          8247 => x"98085482",
          8248 => x"b6980880",
          8249 => x"2eff9b38",
          8250 => x"73842e09",
          8251 => x"81068338",
          8252 => x"87547382",
          8253 => x"b6980c8b",
          8254 => x"3d0d04fd",
          8255 => x"3d0d769a",
          8256 => x"115254eb",
          8257 => x"ec3f82b6",
          8258 => x"980883ff",
          8259 => x"ff067670",
          8260 => x"33515353",
          8261 => x"71832e09",
          8262 => x"81069038",
          8263 => x"941451eb",
          8264 => x"d03f82b6",
          8265 => x"9808902b",
          8266 => x"73075372",
          8267 => x"82b6980c",
          8268 => x"853d0d04",
          8269 => x"fc3d0d77",
          8270 => x"797083ff",
          8271 => x"ff06549a",
          8272 => x"12535555",
          8273 => x"ebed3f76",
          8274 => x"70335153",
          8275 => x"72832e09",
          8276 => x"81068b38",
          8277 => x"73902a52",
          8278 => x"941551eb",
          8279 => x"d63f863d",
          8280 => x"0d04f73d",
          8281 => x"0d7b7d5b",
          8282 => x"55847508",
          8283 => x"5a589815",
          8284 => x"08802e81",
          8285 => x"8a389815",
          8286 => x"08527851",
          8287 => x"ee8f3f82",
          8288 => x"b6980858",
          8289 => x"82b69808",
          8290 => x"80f5389c",
          8291 => x"15087033",
          8292 => x"55537386",
          8293 => x"38845880",
          8294 => x"e6398b13",
          8295 => x"3370bf06",
          8296 => x"7081ff06",
          8297 => x"58515372",
          8298 => x"86163482",
          8299 => x"b6980853",
          8300 => x"7381e52e",
          8301 => x"83388153",
          8302 => x"73ae2ea9",
          8303 => x"38817074",
          8304 => x"06545772",
          8305 => x"802e9e38",
          8306 => x"758f2e99",
          8307 => x"3882b698",
          8308 => x"0876df06",
          8309 => x"54547288",
          8310 => x"2e098106",
          8311 => x"83387654",
          8312 => x"737a2ea0",
          8313 => x"38805274",
          8314 => x"51fafc3f",
          8315 => x"82b69808",
          8316 => x"5882b698",
          8317 => x"08893898",
          8318 => x"1508fefa",
          8319 => x"38863980",
          8320 => x"0b98160c",
          8321 => x"7782b698",
          8322 => x"0c8b3d0d",
          8323 => x"04fb3d0d",
          8324 => x"77700857",
          8325 => x"54815273",
          8326 => x"51fcc53f",
          8327 => x"82b69808",
          8328 => x"5582b698",
          8329 => x"08b43898",
          8330 => x"14085275",
          8331 => x"51ecde3f",
          8332 => x"82b69808",
          8333 => x"5582b698",
          8334 => x"08a038a0",
          8335 => x"5382b698",
          8336 => x"08529c14",
          8337 => x"0851eadb",
          8338 => x"3f8b53a0",
          8339 => x"14529c14",
          8340 => x"0851eaac",
          8341 => x"3f810b83",
          8342 => x"17347482",
          8343 => x"b6980c87",
          8344 => x"3d0d04fd",
          8345 => x"3d0d7570",
          8346 => x"08981208",
          8347 => x"54705355",
          8348 => x"53ec9a3f",
          8349 => x"82b69808",
          8350 => x"8d389c13",
          8351 => x"0853e573",
          8352 => x"34810b83",
          8353 => x"1534853d",
          8354 => x"0d04fa3d",
          8355 => x"0d787a57",
          8356 => x"57800b89",
          8357 => x"17349817",
          8358 => x"08802e81",
          8359 => x"82388070",
          8360 => x"89185555",
          8361 => x"559c1708",
          8362 => x"14703381",
          8363 => x"16565152",
          8364 => x"71a02ea8",
          8365 => x"3871852e",
          8366 => x"09810684",
          8367 => x"3881e552",
          8368 => x"73892e09",
          8369 => x"81068b38",
          8370 => x"ae737081",
          8371 => x"05553481",
          8372 => x"15557173",
          8373 => x"70810555",
          8374 => x"34811555",
          8375 => x"8a7427c5",
          8376 => x"38751588",
          8377 => x"0552800b",
          8378 => x"8113349c",
          8379 => x"1708528b",
          8380 => x"12338817",
          8381 => x"349c1708",
          8382 => x"9c115252",
          8383 => x"e88a3f82",
          8384 => x"b6980876",
          8385 => x"0c961251",
          8386 => x"e7e73f82",
          8387 => x"b6980886",
          8388 => x"17239812",
          8389 => x"51e7da3f",
          8390 => x"82b69808",
          8391 => x"84172388",
          8392 => x"3d0d04f3",
          8393 => x"3d0d7f70",
          8394 => x"085e5b80",
          8395 => x"61703351",
          8396 => x"555573af",
          8397 => x"2e833881",
          8398 => x"557380dc",
          8399 => x"2e913874",
          8400 => x"802e8c38",
          8401 => x"941d0888",
          8402 => x"1c0caa39",
          8403 => x"81154180",
          8404 => x"61703356",
          8405 => x"565673af",
          8406 => x"2e098106",
          8407 => x"83388156",
          8408 => x"7380dc32",
          8409 => x"70307080",
          8410 => x"25780751",
          8411 => x"515473dc",
          8412 => x"3873881c",
          8413 => x"0c607033",
          8414 => x"5154739f",
          8415 => x"269638ff",
          8416 => x"800bab1c",
          8417 => x"3480527a",
          8418 => x"51f6913f",
          8419 => x"82b69808",
          8420 => x"55859839",
          8421 => x"913d61a0",
          8422 => x"1d5c5a5e",
          8423 => x"8b53a052",
          8424 => x"7951e7ff",
          8425 => x"3f807059",
          8426 => x"57887933",
          8427 => x"555c73ae",
          8428 => x"2e098106",
          8429 => x"80d43878",
          8430 => x"18703381",
          8431 => x"1a71ae32",
          8432 => x"7030709f",
          8433 => x"2a738226",
          8434 => x"07515153",
          8435 => x"5a575473",
          8436 => x"8c387917",
          8437 => x"54757434",
          8438 => x"811757db",
          8439 => x"3975af32",
          8440 => x"7030709f",
          8441 => x"2a515154",
          8442 => x"7580dc2e",
          8443 => x"8c387380",
          8444 => x"2e873875",
          8445 => x"a02682bd",
          8446 => x"3877197e",
          8447 => x"0ca454a0",
          8448 => x"762782bd",
          8449 => x"38a05482",
          8450 => x"b8397818",
          8451 => x"7033811a",
          8452 => x"5a5754a0",
          8453 => x"762781fc",
          8454 => x"3875af32",
          8455 => x"70307780",
          8456 => x"dc327030",
          8457 => x"72802571",
          8458 => x"80250751",
          8459 => x"51565155",
          8460 => x"73802eac",
          8461 => x"38843981",
          8462 => x"18588078",
          8463 => x"1a703351",
          8464 => x"555573af",
          8465 => x"2e098106",
          8466 => x"83388155",
          8467 => x"7380dc32",
          8468 => x"70307080",
          8469 => x"25770751",
          8470 => x"515473db",
          8471 => x"3881b539",
          8472 => x"75ae2e09",
          8473 => x"81068338",
          8474 => x"8154767c",
          8475 => x"27740754",
          8476 => x"73802ea2",
          8477 => x"387b8b32",
          8478 => x"703077ae",
          8479 => x"32703072",
          8480 => x"8025719f",
          8481 => x"2a075351",
          8482 => x"56515574",
          8483 => x"81a73888",
          8484 => x"578b5cfe",
          8485 => x"f5397598",
          8486 => x"2b547380",
          8487 => x"258c3875",
          8488 => x"80ff0682",
          8489 => x"afe01133",
          8490 => x"57547551",
          8491 => x"e6e13f82",
          8492 => x"b6980880",
          8493 => x"2eb23878",
          8494 => x"18703381",
          8495 => x"1a71545a",
          8496 => x"5654e6d2",
          8497 => x"3f82b698",
          8498 => x"08802e80",
          8499 => x"e838ff1c",
          8500 => x"54767427",
          8501 => x"80df3879",
          8502 => x"17547574",
          8503 => x"3481177a",
          8504 => x"11555774",
          8505 => x"7434a739",
          8506 => x"755282af",
          8507 => x"8051e5fe",
          8508 => x"3f82b698",
          8509 => x"08bf38ff",
          8510 => x"9f165473",
          8511 => x"99268938",
          8512 => x"e0167081",
          8513 => x"ff065754",
          8514 => x"79175475",
          8515 => x"74348117",
          8516 => x"57fdf739",
          8517 => x"77197e0c",
          8518 => x"76802e99",
          8519 => x"38793354",
          8520 => x"7381e52e",
          8521 => x"09810684",
          8522 => x"38857a34",
          8523 => x"8454a076",
          8524 => x"278f388b",
          8525 => x"39865581",
          8526 => x"f2398456",
          8527 => x"80f33980",
          8528 => x"54738b1b",
          8529 => x"34807b08",
          8530 => x"58527a51",
          8531 => x"f2ce3f82",
          8532 => x"b6980856",
          8533 => x"82b69808",
          8534 => x"80d73898",
          8535 => x"1b085276",
          8536 => x"51e6aa3f",
          8537 => x"82b69808",
          8538 => x"5682b698",
          8539 => x"0880c238",
          8540 => x"9c1b0870",
          8541 => x"33555573",
          8542 => x"802effbe",
          8543 => x"388b1533",
          8544 => x"bf065473",
          8545 => x"861c348b",
          8546 => x"15337083",
          8547 => x"2a708106",
          8548 => x"51555873",
          8549 => x"92388b53",
          8550 => x"79527451",
          8551 => x"e49f3f82",
          8552 => x"b6980880",
          8553 => x"2e8b3875",
          8554 => x"527a51f3",
          8555 => x"ba3fff9f",
          8556 => x"3975ab1c",
          8557 => x"33575574",
          8558 => x"802ebb38",
          8559 => x"74842e09",
          8560 => x"810680e7",
          8561 => x"3875852a",
          8562 => x"70810677",
          8563 => x"822a5851",
          8564 => x"5473802e",
          8565 => x"96387581",
          8566 => x"06547380",
          8567 => x"2efbb538",
          8568 => x"ff800bab",
          8569 => x"1c348055",
          8570 => x"80c13975",
          8571 => x"81065473",
          8572 => x"ba388555",
          8573 => x"b6397582",
          8574 => x"2a708106",
          8575 => x"515473ab",
          8576 => x"38861b33",
          8577 => x"70842a70",
          8578 => x"81065155",
          8579 => x"5573802e",
          8580 => x"e138901b",
          8581 => x"0883ff06",
          8582 => x"1db40552",
          8583 => x"7c51f5db",
          8584 => x"3f82b698",
          8585 => x"08881c0c",
          8586 => x"faea3974",
          8587 => x"82b6980c",
          8588 => x"8f3d0d04",
          8589 => x"f63d0d7c",
          8590 => x"5bff7b08",
          8591 => x"70717355",
          8592 => x"595c5559",
          8593 => x"73802e81",
          8594 => x"c6387570",
          8595 => x"81055733",
          8596 => x"70a02652",
          8597 => x"5271ba2e",
          8598 => x"8d3870ee",
          8599 => x"3871ba2e",
          8600 => x"09810681",
          8601 => x"a5387333",
          8602 => x"d0117081",
          8603 => x"ff065152",
          8604 => x"53708926",
          8605 => x"91388214",
          8606 => x"7381ff06",
          8607 => x"d0055652",
          8608 => x"71762e80",
          8609 => x"f738800b",
          8610 => x"82afd059",
          8611 => x"5577087a",
          8612 => x"55577670",
          8613 => x"81055833",
          8614 => x"74708105",
          8615 => x"5633ff9f",
          8616 => x"12535353",
          8617 => x"70992689",
          8618 => x"38e01370",
          8619 => x"81ff0654",
          8620 => x"51ff9f12",
          8621 => x"51709926",
          8622 => x"8938e012",
          8623 => x"7081ff06",
          8624 => x"53517230",
          8625 => x"709f2a51",
          8626 => x"5172722e",
          8627 => x"09810685",
          8628 => x"3870ffbe",
          8629 => x"38723074",
          8630 => x"77327030",
          8631 => x"7072079f",
          8632 => x"2a739f2a",
          8633 => x"07535454",
          8634 => x"5170802e",
          8635 => x"8f388115",
          8636 => x"84195955",
          8637 => x"837525ff",
          8638 => x"94388b39",
          8639 => x"74832486",
          8640 => x"3874767c",
          8641 => x"0c597851",
          8642 => x"863982cd",
          8643 => x"e4335170",
          8644 => x"82b6980c",
          8645 => x"8c3d0d04",
          8646 => x"fa3d0d78",
          8647 => x"56800b83",
          8648 => x"1734ff0b",
          8649 => x"b0170c79",
          8650 => x"527551e2",
          8651 => x"e03f8455",
          8652 => x"82b69808",
          8653 => x"81803884",
          8654 => x"b21651df",
          8655 => x"b43f82b6",
          8656 => x"980883ff",
          8657 => x"ff065483",
          8658 => x"557382d4",
          8659 => x"d52e0981",
          8660 => x"0680e338",
          8661 => x"800bb417",
          8662 => x"33565774",
          8663 => x"81e92e09",
          8664 => x"81068338",
          8665 => x"81577481",
          8666 => x"eb327030",
          8667 => x"70802579",
          8668 => x"07515154",
          8669 => x"738a3874",
          8670 => x"81e82e09",
          8671 => x"8106b538",
          8672 => x"835382af",
          8673 => x"905280ea",
          8674 => x"1651e0b1",
          8675 => x"3f82b698",
          8676 => x"085582b6",
          8677 => x"9808802e",
          8678 => x"9d388553",
          8679 => x"82af9452",
          8680 => x"81861651",
          8681 => x"e0973f82",
          8682 => x"b6980855",
          8683 => x"82b69808",
          8684 => x"802e8338",
          8685 => x"82557482",
          8686 => x"b6980c88",
          8687 => x"3d0d04f2",
          8688 => x"3d0d6102",
          8689 => x"840580cb",
          8690 => x"05335855",
          8691 => x"80750c60",
          8692 => x"51fce13f",
          8693 => x"82b69808",
          8694 => x"588b5680",
          8695 => x"0b82b698",
          8696 => x"082486fc",
          8697 => x"3882b698",
          8698 => x"08842982",
          8699 => x"cdd00570",
          8700 => x"0855538c",
          8701 => x"5673802e",
          8702 => x"86e63873",
          8703 => x"750c7681",
          8704 => x"fe067433",
          8705 => x"54577280",
          8706 => x"2eae3881",
          8707 => x"143351d7",
          8708 => x"ca3f82b6",
          8709 => x"980881ff",
          8710 => x"06708106",
          8711 => x"54557298",
          8712 => x"3876802e",
          8713 => x"86b83874",
          8714 => x"822a7081",
          8715 => x"0651538a",
          8716 => x"567286ac",
          8717 => x"3886a739",
          8718 => x"80743477",
          8719 => x"81153481",
          8720 => x"52811433",
          8721 => x"51d7b23f",
          8722 => x"82b69808",
          8723 => x"81ff0670",
          8724 => x"81065455",
          8725 => x"83567286",
          8726 => x"87387680",
          8727 => x"2e8f3874",
          8728 => x"822a7081",
          8729 => x"0651538a",
          8730 => x"567285f4",
          8731 => x"38807053",
          8732 => x"74525bfd",
          8733 => x"a33f82b6",
          8734 => x"980881ff",
          8735 => x"06577682",
          8736 => x"2e098106",
          8737 => x"80e2388c",
          8738 => x"3d745658",
          8739 => x"835683f6",
          8740 => x"15337058",
          8741 => x"5372802e",
          8742 => x"8d3883fa",
          8743 => x"1551dce8",
          8744 => x"3f82b698",
          8745 => x"08577678",
          8746 => x"7084055a",
          8747 => x"0cff1690",
          8748 => x"16565675",
          8749 => x"8025d738",
          8750 => x"800b8d3d",
          8751 => x"54567270",
          8752 => x"84055408",
          8753 => x"5b83577a",
          8754 => x"802e9538",
          8755 => x"7a527351",
          8756 => x"fcc63f82",
          8757 => x"b6980881",
          8758 => x"ff065781",
          8759 => x"77278938",
          8760 => x"81165683",
          8761 => x"7627d738",
          8762 => x"81567684",
          8763 => x"2e84f138",
          8764 => x"8d567681",
          8765 => x"2684e938",
          8766 => x"bf1451db",
          8767 => x"f43f82b6",
          8768 => x"980883ff",
          8769 => x"ff065372",
          8770 => x"84802e09",
          8771 => x"810684d0",
          8772 => x"3880ca14",
          8773 => x"51dbda3f",
          8774 => x"82b69808",
          8775 => x"83ffff06",
          8776 => x"58778d38",
          8777 => x"80d81451",
          8778 => x"dbde3f82",
          8779 => x"b6980858",
          8780 => x"779c150c",
          8781 => x"80c41433",
          8782 => x"82153480",
          8783 => x"c41433ff",
          8784 => x"117081ff",
          8785 => x"06515455",
          8786 => x"8d567281",
          8787 => x"26849138",
          8788 => x"7481ff06",
          8789 => x"78712980",
          8790 => x"c1163352",
          8791 => x"5953728a",
          8792 => x"15237280",
          8793 => x"2e8b38ff",
          8794 => x"13730653",
          8795 => x"72802e86",
          8796 => x"388d5683",
          8797 => x"eb3980c5",
          8798 => x"1451daf5",
          8799 => x"3f82b698",
          8800 => x"085382b6",
          8801 => x"98088815",
          8802 => x"23728f06",
          8803 => x"578d5676",
          8804 => x"83ce3880",
          8805 => x"c71451da",
          8806 => x"d83f82b6",
          8807 => x"980883ff",
          8808 => x"ff065574",
          8809 => x"8d3880d4",
          8810 => x"1451dadc",
          8811 => x"3f82b698",
          8812 => x"085580c2",
          8813 => x"1451dab9",
          8814 => x"3f82b698",
          8815 => x"0883ffff",
          8816 => x"06538d56",
          8817 => x"72802e83",
          8818 => x"97388814",
          8819 => x"22781471",
          8820 => x"842a055a",
          8821 => x"5a787526",
          8822 => x"8386388a",
          8823 => x"14225274",
          8824 => x"793151fe",
          8825 => x"f39d3f82",
          8826 => x"b6980855",
          8827 => x"82b69808",
          8828 => x"802e82ec",
          8829 => x"3882b698",
          8830 => x"0880ffff",
          8831 => x"fff52683",
          8832 => x"38835774",
          8833 => x"83fff526",
          8834 => x"83388257",
          8835 => x"749ff526",
          8836 => x"85388157",
          8837 => x"89398d56",
          8838 => x"76802e82",
          8839 => x"c3388215",
          8840 => x"7098160c",
          8841 => x"7ba0160c",
          8842 => x"731c70a4",
          8843 => x"170c7a1d",
          8844 => x"ac170c54",
          8845 => x"5576832e",
          8846 => x"098106af",
          8847 => x"3880de14",
          8848 => x"51d9ae3f",
          8849 => x"82b69808",
          8850 => x"83ffff06",
          8851 => x"538d5672",
          8852 => x"828e3879",
          8853 => x"828a3880",
          8854 => x"e01451d9",
          8855 => x"ab3f82b6",
          8856 => x"9808a815",
          8857 => x"0c74822b",
          8858 => x"53a2398d",
          8859 => x"5679802e",
          8860 => x"81ee3877",
          8861 => x"13a8150c",
          8862 => x"74155376",
          8863 => x"822e8d38",
          8864 => x"74101570",
          8865 => x"812a7681",
          8866 => x"06055153",
          8867 => x"83ff1389",
          8868 => x"2a538d56",
          8869 => x"729c1508",
          8870 => x"2681c538",
          8871 => x"ff0b9015",
          8872 => x"0cff0b8c",
          8873 => x"150cff80",
          8874 => x"0b841534",
          8875 => x"76832e09",
          8876 => x"81068192",
          8877 => x"3880e414",
          8878 => x"51d8b63f",
          8879 => x"82b69808",
          8880 => x"83ffff06",
          8881 => x"5372812e",
          8882 => x"09810680",
          8883 => x"f938811b",
          8884 => x"527351db",
          8885 => x"b83f82b6",
          8886 => x"980880ea",
          8887 => x"3882b698",
          8888 => x"08841534",
          8889 => x"84b21451",
          8890 => x"d8873f82",
          8891 => x"b6980883",
          8892 => x"ffff0653",
          8893 => x"7282d4d5",
          8894 => x"2e098106",
          8895 => x"80c838b4",
          8896 => x"1451d884",
          8897 => x"3f82b698",
          8898 => x"08848b85",
          8899 => x"a4d22e09",
          8900 => x"8106b338",
          8901 => x"84981451",
          8902 => x"d7ee3f82",
          8903 => x"b6980886",
          8904 => x"8a85e4f2",
          8905 => x"2e098106",
          8906 => x"9d38849c",
          8907 => x"1451d7d8",
          8908 => x"3f82b698",
          8909 => x"0890150c",
          8910 => x"84a01451",
          8911 => x"d7ca3f82",
          8912 => x"b698088c",
          8913 => x"150c7674",
          8914 => x"3482cde0",
          8915 => x"22810553",
          8916 => x"7282cde0",
          8917 => x"23728615",
          8918 => x"23800b94",
          8919 => x"150c8056",
          8920 => x"7582b698",
          8921 => x"0c903d0d",
          8922 => x"04fb3d0d",
          8923 => x"77548955",
          8924 => x"73802eb9",
          8925 => x"38730853",
          8926 => x"72802eb1",
          8927 => x"38723352",
          8928 => x"71802ea9",
          8929 => x"38861322",
          8930 => x"84152257",
          8931 => x"5271762e",
          8932 => x"09810699",
          8933 => x"38811333",
          8934 => x"51d0c03f",
          8935 => x"82b69808",
          8936 => x"81065271",
          8937 => x"88387174",
          8938 => x"08545583",
          8939 => x"39805378",
          8940 => x"73710c52",
          8941 => x"7482b698",
          8942 => x"0c873d0d",
          8943 => x"04fa3d0d",
          8944 => x"02ab0533",
          8945 => x"7a58893d",
          8946 => x"fc055256",
          8947 => x"f4e63f8b",
          8948 => x"54800b82",
          8949 => x"b6980824",
          8950 => x"bc3882b6",
          8951 => x"98088429",
          8952 => x"82cdd005",
          8953 => x"70085555",
          8954 => x"73802e84",
          8955 => x"38807434",
          8956 => x"78547380",
          8957 => x"2e843880",
          8958 => x"74347875",
          8959 => x"0c755475",
          8960 => x"802e9238",
          8961 => x"8053893d",
          8962 => x"70538405",
          8963 => x"51f7b03f",
          8964 => x"82b69808",
          8965 => x"547382b6",
          8966 => x"980c883d",
          8967 => x"0d04eb3d",
          8968 => x"0d670284",
          8969 => x"0580e705",
          8970 => x"33595989",
          8971 => x"5478802e",
          8972 => x"84c83877",
          8973 => x"bf067054",
          8974 => x"983dd005",
          8975 => x"53993d84",
          8976 => x"055258f6",
          8977 => x"fa3f82b6",
          8978 => x"98085582",
          8979 => x"b6980884",
          8980 => x"a4387a5c",
          8981 => x"68528c3d",
          8982 => x"705256ed",
          8983 => x"c63f82b6",
          8984 => x"98085582",
          8985 => x"b6980892",
          8986 => x"380280d7",
          8987 => x"05337098",
          8988 => x"2b555773",
          8989 => x"80258338",
          8990 => x"8655779c",
          8991 => x"06547380",
          8992 => x"2e81ab38",
          8993 => x"74802e95",
          8994 => x"3874842e",
          8995 => x"098106aa",
          8996 => x"387551ea",
          8997 => x"f83f82b6",
          8998 => x"9808559e",
          8999 => x"3902b205",
          9000 => x"33910654",
          9001 => x"7381b838",
          9002 => x"77822a70",
          9003 => x"81065154",
          9004 => x"73802e8e",
          9005 => x"38885583",
          9006 => x"bc397788",
          9007 => x"07587483",
          9008 => x"b4387783",
          9009 => x"2a708106",
          9010 => x"51547380",
          9011 => x"2e81af38",
          9012 => x"62527a51",
          9013 => x"e8a53f82",
          9014 => x"b6980856",
          9015 => x"8288b20a",
          9016 => x"52628e05",
          9017 => x"51d4ea3f",
          9018 => x"6254a00b",
          9019 => x"8b153480",
          9020 => x"5362527a",
          9021 => x"51e8bd3f",
          9022 => x"8052629c",
          9023 => x"0551d4d1",
          9024 => x"3f7a5481",
          9025 => x"0b831534",
          9026 => x"75802e80",
          9027 => x"f1387ab0",
          9028 => x"11085154",
          9029 => x"80537552",
          9030 => x"973dd405",
          9031 => x"51ddbe3f",
          9032 => x"82b69808",
          9033 => x"5582b698",
          9034 => x"0882ca38",
          9035 => x"b7397482",
          9036 => x"c43802b2",
          9037 => x"05337084",
          9038 => x"2a708106",
          9039 => x"51555673",
          9040 => x"802e8638",
          9041 => x"845582ad",
          9042 => x"3977812a",
          9043 => x"70810651",
          9044 => x"5473802e",
          9045 => x"a9387581",
          9046 => x"06547380",
          9047 => x"2ea03887",
          9048 => x"55829239",
          9049 => x"73527a51",
          9050 => x"d6a33f82",
          9051 => x"b698087b",
          9052 => x"ff188c12",
          9053 => x"0c555582",
          9054 => x"b6980881",
          9055 => x"f8387783",
          9056 => x"2a708106",
          9057 => x"51547380",
          9058 => x"2e863877",
          9059 => x"80c00758",
          9060 => x"7ab01108",
          9061 => x"a01b0c63",
          9062 => x"a41b0c63",
          9063 => x"53705257",
          9064 => x"e6d93f82",
          9065 => x"b6980882",
          9066 => x"b6980888",
          9067 => x"1b0c639c",
          9068 => x"05525ad2",
          9069 => x"d33f82b6",
          9070 => x"980882b6",
          9071 => x"98088c1b",
          9072 => x"0c777a0c",
          9073 => x"56861722",
          9074 => x"841a2377",
          9075 => x"901a3480",
          9076 => x"0b911a34",
          9077 => x"800b9c1a",
          9078 => x"0c800b94",
          9079 => x"1a0c7785",
          9080 => x"2a708106",
          9081 => x"51547380",
          9082 => x"2e818d38",
          9083 => x"82b69808",
          9084 => x"802e8184",
          9085 => x"3882b698",
          9086 => x"08941a0c",
          9087 => x"8a172270",
          9088 => x"892b7b52",
          9089 => x"5957a839",
          9090 => x"76527851",
          9091 => x"d79f3f82",
          9092 => x"b6980857",
          9093 => x"82b69808",
          9094 => x"81268338",
          9095 => x"825582b6",
          9096 => x"9808ff2e",
          9097 => x"09810683",
          9098 => x"38795575",
          9099 => x"78315674",
          9100 => x"30707607",
          9101 => x"80255154",
          9102 => x"7776278a",
          9103 => x"38817075",
          9104 => x"06555a73",
          9105 => x"c3387698",
          9106 => x"1a0c74a9",
          9107 => x"387583ff",
          9108 => x"06547380",
          9109 => x"2ea23876",
          9110 => x"527a51d6",
          9111 => x"a63f82b6",
          9112 => x"98088538",
          9113 => x"82558e39",
          9114 => x"75892a82",
          9115 => x"b6980805",
          9116 => x"9c1a0c84",
          9117 => x"3980790c",
          9118 => x"74547382",
          9119 => x"b6980c97",
          9120 => x"3d0d04f2",
          9121 => x"3d0d6063",
          9122 => x"65644040",
          9123 => x"5d59807e",
          9124 => x"0c903dfc",
          9125 => x"05527851",
          9126 => x"f9cf3f82",
          9127 => x"b6980855",
          9128 => x"82b69808",
          9129 => x"8a389119",
          9130 => x"33557480",
          9131 => x"2e863874",
          9132 => x"5682c439",
          9133 => x"90193381",
          9134 => x"06558756",
          9135 => x"74802e82",
          9136 => x"b6389539",
          9137 => x"820b911a",
          9138 => x"34825682",
          9139 => x"aa39810b",
          9140 => x"911a3481",
          9141 => x"5682a039",
          9142 => x"8c190894",
          9143 => x"1a083155",
          9144 => x"747c2783",
          9145 => x"38745c7b",
          9146 => x"802e8289",
          9147 => x"38941908",
          9148 => x"7083ff06",
          9149 => x"56567481",
          9150 => x"b2387e8a",
          9151 => x"1122ff05",
          9152 => x"77892a06",
          9153 => x"5b5579a8",
          9154 => x"38758738",
          9155 => x"88190855",
          9156 => x"8f399819",
          9157 => x"08527851",
          9158 => x"d5933f82",
          9159 => x"b6980855",
          9160 => x"817527ff",
          9161 => x"9f3874ff",
          9162 => x"2effa338",
          9163 => x"74981a0c",
          9164 => x"98190852",
          9165 => x"7e51d4cb",
          9166 => x"3f82b698",
          9167 => x"08802eff",
          9168 => x"833882b6",
          9169 => x"98081a7c",
          9170 => x"892a5957",
          9171 => x"77802e80",
          9172 => x"d638771a",
          9173 => x"7f8a1122",
          9174 => x"585c5575",
          9175 => x"75278538",
          9176 => x"757a3158",
          9177 => x"77547653",
          9178 => x"7c52811b",
          9179 => x"3351ca88",
          9180 => x"3f82b698",
          9181 => x"08fed738",
          9182 => x"7e831133",
          9183 => x"56567480",
          9184 => x"2e9f38b0",
          9185 => x"16087731",
          9186 => x"55747827",
          9187 => x"94388480",
          9188 => x"53b41652",
          9189 => x"b0160877",
          9190 => x"31892b7d",
          9191 => x"0551cfe0",
          9192 => x"3f77892b",
          9193 => x"56b93976",
          9194 => x"9c1a0c94",
          9195 => x"190883ff",
          9196 => x"06848071",
          9197 => x"3157557b",
          9198 => x"76278338",
          9199 => x"7b569c19",
          9200 => x"08527e51",
          9201 => x"d1c73f82",
          9202 => x"b69808fe",
          9203 => x"81387553",
          9204 => x"94190883",
          9205 => x"ff061fb4",
          9206 => x"05527c51",
          9207 => x"cfa23f7b",
          9208 => x"76317e08",
          9209 => x"177f0c76",
          9210 => x"1e941b08",
          9211 => x"18941c0c",
          9212 => x"5e5cfdf3",
          9213 => x"39805675",
          9214 => x"82b6980c",
          9215 => x"903d0d04",
          9216 => x"f23d0d60",
          9217 => x"63656440",
          9218 => x"405d5880",
          9219 => x"7e0c903d",
          9220 => x"fc055277",
          9221 => x"51f6d23f",
          9222 => x"82b69808",
          9223 => x"5582b698",
          9224 => x"088a3891",
          9225 => x"18335574",
          9226 => x"802e8638",
          9227 => x"745683b8",
          9228 => x"39901833",
          9229 => x"70812a70",
          9230 => x"81065156",
          9231 => x"56875674",
          9232 => x"802e83a4",
          9233 => x"38953982",
          9234 => x"0b911934",
          9235 => x"82568398",
          9236 => x"39810b91",
          9237 => x"19348156",
          9238 => x"838e3994",
          9239 => x"18087c11",
          9240 => x"56567476",
          9241 => x"27843875",
          9242 => x"095c7b80",
          9243 => x"2e82ec38",
          9244 => x"94180870",
          9245 => x"83ff0656",
          9246 => x"567481fd",
          9247 => x"387e8a11",
          9248 => x"22ff0577",
          9249 => x"892a065c",
          9250 => x"557abf38",
          9251 => x"758c3888",
          9252 => x"18085574",
          9253 => x"9c387a52",
          9254 => x"85399818",
          9255 => x"08527751",
          9256 => x"d7e73f82",
          9257 => x"b6980855",
          9258 => x"82b69808",
          9259 => x"802e82ab",
          9260 => x"3874812e",
          9261 => x"ff913874",
          9262 => x"ff2eff95",
          9263 => x"38749819",
          9264 => x"0c881808",
          9265 => x"85387488",
          9266 => x"190c7e55",
          9267 => x"b015089c",
          9268 => x"19082e09",
          9269 => x"81068d38",
          9270 => x"7451cec1",
          9271 => x"3f82b698",
          9272 => x"08feee38",
          9273 => x"98180852",
          9274 => x"7e51d197",
          9275 => x"3f82b698",
          9276 => x"08802efe",
          9277 => x"d23882b6",
          9278 => x"98081b7c",
          9279 => x"892a5a57",
          9280 => x"78802e80",
          9281 => x"d538781b",
          9282 => x"7f8a1122",
          9283 => x"585b5575",
          9284 => x"75278538",
          9285 => x"757b3159",
          9286 => x"78547653",
          9287 => x"7c52811a",
          9288 => x"3351c8be",
          9289 => x"3f82b698",
          9290 => x"08fea638",
          9291 => x"7eb01108",
          9292 => x"78315656",
          9293 => x"7479279b",
          9294 => x"38848053",
          9295 => x"b0160877",
          9296 => x"31892b7d",
          9297 => x"0552b416",
          9298 => x"51ccb53f",
          9299 => x"7e55800b",
          9300 => x"83163478",
          9301 => x"892b5680",
          9302 => x"db398c18",
          9303 => x"08941908",
          9304 => x"2693387e",
          9305 => x"51cdb63f",
          9306 => x"82b69808",
          9307 => x"fde3387e",
          9308 => x"77b0120c",
          9309 => x"55769c19",
          9310 => x"0c941808",
          9311 => x"83ff0684",
          9312 => x"80713157",
          9313 => x"557b7627",
          9314 => x"83387b56",
          9315 => x"9c180852",
          9316 => x"7e51cdf9",
          9317 => x"3f82b698",
          9318 => x"08fdb638",
          9319 => x"75537c52",
          9320 => x"94180883",
          9321 => x"ff061fb4",
          9322 => x"0551cbd4",
          9323 => x"3f7e5581",
          9324 => x"0b831634",
          9325 => x"7b76317e",
          9326 => x"08177f0c",
          9327 => x"761e941a",
          9328 => x"08187094",
          9329 => x"1c0c8c1b",
          9330 => x"0858585e",
          9331 => x"5c747627",
          9332 => x"83387555",
          9333 => x"748c190c",
          9334 => x"fd903990",
          9335 => x"183380c0",
          9336 => x"07557490",
          9337 => x"19348056",
          9338 => x"7582b698",
          9339 => x"0c903d0d",
          9340 => x"04f83d0d",
          9341 => x"7a8b3dfc",
          9342 => x"05537052",
          9343 => x"56f2ea3f",
          9344 => x"82b69808",
          9345 => x"5782b698",
          9346 => x"0880fb38",
          9347 => x"90163370",
          9348 => x"862a7081",
          9349 => x"06515555",
          9350 => x"73802e80",
          9351 => x"e938a016",
          9352 => x"08527851",
          9353 => x"cce73f82",
          9354 => x"b6980857",
          9355 => x"82b69808",
          9356 => x"80d438a4",
          9357 => x"16088b11",
          9358 => x"33a00755",
          9359 => x"55738b16",
          9360 => x"34881608",
          9361 => x"53745275",
          9362 => x"0851dde8",
          9363 => x"3f8c1608",
          9364 => x"529c1551",
          9365 => x"c9fb3f82",
          9366 => x"88b20a52",
          9367 => x"961551c9",
          9368 => x"f03f7652",
          9369 => x"921551c9",
          9370 => x"ca3f7854",
          9371 => x"810b8315",
          9372 => x"347851cc",
          9373 => x"df3f82b6",
          9374 => x"98089017",
          9375 => x"3381bf06",
          9376 => x"55577390",
          9377 => x"17347682",
          9378 => x"b6980c8a",
          9379 => x"3d0d04fc",
          9380 => x"3d0d7670",
          9381 => x"5254fed9",
          9382 => x"3f82b698",
          9383 => x"085382b6",
          9384 => x"98089c38",
          9385 => x"863dfc05",
          9386 => x"527351f1",
          9387 => x"bc3f82b6",
          9388 => x"98085382",
          9389 => x"b6980887",
          9390 => x"3882b698",
          9391 => x"08740c72",
          9392 => x"82b6980c",
          9393 => x"863d0d04",
          9394 => x"ff3d0d84",
          9395 => x"3d51e6e4",
          9396 => x"3f8b5280",
          9397 => x"0b82b698",
          9398 => x"08248b38",
          9399 => x"82b69808",
          9400 => x"82cde434",
          9401 => x"80527182",
          9402 => x"b6980c83",
          9403 => x"3d0d04ef",
          9404 => x"3d0d8053",
          9405 => x"933dd005",
          9406 => x"52943d51",
          9407 => x"e9c13f82",
          9408 => x"b6980855",
          9409 => x"82b69808",
          9410 => x"80e03876",
          9411 => x"58635293",
          9412 => x"3dd40551",
          9413 => x"e08d3f82",
          9414 => x"b6980855",
          9415 => x"82b69808",
          9416 => x"bc380280",
          9417 => x"c7053370",
          9418 => x"982b5556",
          9419 => x"73802589",
          9420 => x"38767a94",
          9421 => x"120c54b2",
          9422 => x"3902a205",
          9423 => x"3370842a",
          9424 => x"70810651",
          9425 => x"55567380",
          9426 => x"2e9e3876",
          9427 => x"7f537052",
          9428 => x"54dba83f",
          9429 => x"82b69808",
          9430 => x"94150c8e",
          9431 => x"3982b698",
          9432 => x"08842e09",
          9433 => x"81068338",
          9434 => x"85557482",
          9435 => x"b6980c93",
          9436 => x"3d0d04e4",
          9437 => x"3d0d6f6f",
          9438 => x"5b5b807a",
          9439 => x"3480539e",
          9440 => x"3dffb805",
          9441 => x"529f3d51",
          9442 => x"e8b53f82",
          9443 => x"b6980857",
          9444 => x"82b69808",
          9445 => x"82fc387b",
          9446 => x"437a7c94",
          9447 => x"11084755",
          9448 => x"58645473",
          9449 => x"802e81ed",
          9450 => x"38a05293",
          9451 => x"3d705255",
          9452 => x"d5ea3f82",
          9453 => x"b6980857",
          9454 => x"82b69808",
          9455 => x"82d43868",
          9456 => x"527b51c9",
          9457 => x"c83f82b6",
          9458 => x"98085782",
          9459 => x"b6980882",
          9460 => x"c1386952",
          9461 => x"7b51daa3",
          9462 => x"3f82b698",
          9463 => x"08457652",
          9464 => x"7451d5b8",
          9465 => x"3f82b698",
          9466 => x"085782b6",
          9467 => x"980882a2",
          9468 => x"38805274",
          9469 => x"51daeb3f",
          9470 => x"82b69808",
          9471 => x"5782b698",
          9472 => x"08a43869",
          9473 => x"527b51d9",
          9474 => x"f23f7382",
          9475 => x"b698082e",
          9476 => x"a6387652",
          9477 => x"7451d6cf",
          9478 => x"3f82b698",
          9479 => x"085782b6",
          9480 => x"9808802e",
          9481 => x"cc387684",
          9482 => x"2e098106",
          9483 => x"86388257",
          9484 => x"81e03976",
          9485 => x"81dc389e",
          9486 => x"3dffbc05",
          9487 => x"527451dc",
          9488 => x"c93f7690",
          9489 => x"3d781181",
          9490 => x"11335156",
          9491 => x"5a567380",
          9492 => x"2e913802",
          9493 => x"b9055581",
          9494 => x"16811670",
          9495 => x"33565656",
          9496 => x"73f53881",
          9497 => x"16547378",
          9498 => x"26819038",
          9499 => x"75802e99",
          9500 => x"38781681",
          9501 => x"0555ff18",
          9502 => x"6f11ff18",
          9503 => x"ff185858",
          9504 => x"55587433",
          9505 => x"743475ee",
          9506 => x"38ff186f",
          9507 => x"115558af",
          9508 => x"7434fe8d",
          9509 => x"39777b2e",
          9510 => x"0981068a",
          9511 => x"38ff186f",
          9512 => x"115558af",
          9513 => x"7434800b",
          9514 => x"82cde433",
          9515 => x"70842982",
          9516 => x"afd00570",
          9517 => x"08703352",
          9518 => x"5c565656",
          9519 => x"73762e8d",
          9520 => x"38811670",
          9521 => x"1a703351",
          9522 => x"555673f5",
          9523 => x"38821654",
          9524 => x"737826a7",
          9525 => x"38805574",
          9526 => x"76279138",
          9527 => x"74195473",
          9528 => x"337a7081",
          9529 => x"055c3481",
          9530 => x"1555ec39",
          9531 => x"ba7a7081",
          9532 => x"055c3474",
          9533 => x"ff2e0981",
          9534 => x"06853891",
          9535 => x"5794396e",
          9536 => x"18811959",
          9537 => x"5473337a",
          9538 => x"7081055c",
          9539 => x"347a7826",
          9540 => x"ee38807a",
          9541 => x"347682b6",
          9542 => x"980c9e3d",
          9543 => x"0d04f73d",
          9544 => x"0d7b7d8d",
          9545 => x"3dfc0554",
          9546 => x"71535755",
          9547 => x"ecbb3f82",
          9548 => x"b6980853",
          9549 => x"82b69808",
          9550 => x"82fa3891",
          9551 => x"15335372",
          9552 => x"82f2388c",
          9553 => x"15085473",
          9554 => x"76279238",
          9555 => x"90153370",
          9556 => x"812a7081",
          9557 => x"06515457",
          9558 => x"72833873",
          9559 => x"56941508",
          9560 => x"54807094",
          9561 => x"170c5875",
          9562 => x"782e8297",
          9563 => x"38798a11",
          9564 => x"2270892b",
          9565 => x"59515373",
          9566 => x"782eb738",
          9567 => x"7652ff16",
          9568 => x"51fedbff",
          9569 => x"3f82b698",
          9570 => x"08ff1578",
          9571 => x"54705355",
          9572 => x"53fedbef",
          9573 => x"3f82b698",
          9574 => x"08732696",
          9575 => x"38763070",
          9576 => x"75067094",
          9577 => x"180c7771",
          9578 => x"31981808",
          9579 => x"57585153",
          9580 => x"b1398815",
          9581 => x"085473a6",
          9582 => x"38735274",
          9583 => x"51cdca3f",
          9584 => x"82b69808",
          9585 => x"5482b698",
          9586 => x"08812e81",
          9587 => x"9a3882b6",
          9588 => x"9808ff2e",
          9589 => x"819b3882",
          9590 => x"b6980888",
          9591 => x"160c7398",
          9592 => x"160c7380",
          9593 => x"2e819c38",
          9594 => x"76762780",
          9595 => x"dc387577",
          9596 => x"31941608",
          9597 => x"1894170c",
          9598 => x"90163370",
          9599 => x"812a7081",
          9600 => x"0651555a",
          9601 => x"5672802e",
          9602 => x"9a387352",
          9603 => x"7451ccf9",
          9604 => x"3f82b698",
          9605 => x"085482b6",
          9606 => x"98089438",
          9607 => x"82b69808",
          9608 => x"56a73973",
          9609 => x"527451c7",
          9610 => x"843f82b6",
          9611 => x"98085473",
          9612 => x"ff2ebe38",
          9613 => x"817427af",
          9614 => x"38795373",
          9615 => x"98140827",
          9616 => x"a6387398",
          9617 => x"160cffa0",
          9618 => x"39941508",
          9619 => x"1694160c",
          9620 => x"7583ff06",
          9621 => x"5372802e",
          9622 => x"aa387352",
          9623 => x"7951c6a3",
          9624 => x"3f82b698",
          9625 => x"08943882",
          9626 => x"0b911634",
          9627 => x"825380c4",
          9628 => x"39810b91",
          9629 => x"16348153",
          9630 => x"bb397589",
          9631 => x"2a82b698",
          9632 => x"08055894",
          9633 => x"1508548c",
          9634 => x"15087427",
          9635 => x"9038738c",
          9636 => x"160c9015",
          9637 => x"3380c007",
          9638 => x"53729016",
          9639 => x"347383ff",
          9640 => x"06537280",
          9641 => x"2e8c3877",
          9642 => x"9c16082e",
          9643 => x"8538779c",
          9644 => x"160c8053",
          9645 => x"7282b698",
          9646 => x"0c8b3d0d",
          9647 => x"04f93d0d",
          9648 => x"79568954",
          9649 => x"75802e81",
          9650 => x"8a388053",
          9651 => x"893dfc05",
          9652 => x"528a3d84",
          9653 => x"0551e1e7",
          9654 => x"3f82b698",
          9655 => x"085582b6",
          9656 => x"980880ea",
          9657 => x"3877760c",
          9658 => x"7a527551",
          9659 => x"d8b53f82",
          9660 => x"b6980855",
          9661 => x"82b69808",
          9662 => x"80c338ab",
          9663 => x"16337098",
          9664 => x"2b555780",
          9665 => x"7424a238",
          9666 => x"86163370",
          9667 => x"842a7081",
          9668 => x"06515557",
          9669 => x"73802ead",
          9670 => x"389c1608",
          9671 => x"527751d3",
          9672 => x"da3f82b6",
          9673 => x"98088817",
          9674 => x"0c775486",
          9675 => x"14228417",
          9676 => x"23745275",
          9677 => x"51cee53f",
          9678 => x"82b69808",
          9679 => x"5574842e",
          9680 => x"09810685",
          9681 => x"38855586",
          9682 => x"3974802e",
          9683 => x"84388076",
          9684 => x"0c745473",
          9685 => x"82b6980c",
          9686 => x"893d0d04",
          9687 => x"fc3d0d76",
          9688 => x"873dfc05",
          9689 => x"53705253",
          9690 => x"e7ff3f82",
          9691 => x"b6980887",
          9692 => x"3882b698",
          9693 => x"08730c86",
          9694 => x"3d0d04fb",
          9695 => x"3d0d7779",
          9696 => x"893dfc05",
          9697 => x"54715356",
          9698 => x"54e7de3f",
          9699 => x"82b69808",
          9700 => x"5382b698",
          9701 => x"0880df38",
          9702 => x"74933882",
          9703 => x"b6980852",
          9704 => x"7351cdf8",
          9705 => x"3f82b698",
          9706 => x"085380ca",
          9707 => x"3982b698",
          9708 => x"08527351",
          9709 => x"d3ac3f82",
          9710 => x"b6980853",
          9711 => x"82b69808",
          9712 => x"842e0981",
          9713 => x"06853880",
          9714 => x"53873982",
          9715 => x"b69808a6",
          9716 => x"38745273",
          9717 => x"51d5b33f",
          9718 => x"72527351",
          9719 => x"cf893f82",
          9720 => x"b6980884",
          9721 => x"32703070",
          9722 => x"72079f2c",
          9723 => x"7082b698",
          9724 => x"08065151",
          9725 => x"54547282",
          9726 => x"b6980c87",
          9727 => x"3d0d04ee",
          9728 => x"3d0d6557",
          9729 => x"8053893d",
          9730 => x"7053963d",
          9731 => x"5256dfaf",
          9732 => x"3f82b698",
          9733 => x"085582b6",
          9734 => x"9808b238",
          9735 => x"64527551",
          9736 => x"d6813f82",
          9737 => x"b6980855",
          9738 => x"82b69808",
          9739 => x"a0380280",
          9740 => x"cb053370",
          9741 => x"982b5558",
          9742 => x"73802585",
          9743 => x"3886558d",
          9744 => x"3976802e",
          9745 => x"88387652",
          9746 => x"7551d4be",
          9747 => x"3f7482b6",
          9748 => x"980c943d",
          9749 => x"0d04f03d",
          9750 => x"0d636555",
          9751 => x"5c805392",
          9752 => x"3dec0552",
          9753 => x"933d51de",
          9754 => x"d63f82b6",
          9755 => x"98085b82",
          9756 => x"b6980882",
          9757 => x"80387c74",
          9758 => x"0c730898",
          9759 => x"1108fe11",
          9760 => x"90130859",
          9761 => x"56585575",
          9762 => x"74269138",
          9763 => x"757c0c81",
          9764 => x"e439815b",
          9765 => x"81cc3982",
          9766 => x"5b81c739",
          9767 => x"82b69808",
          9768 => x"75335559",
          9769 => x"73812e09",
          9770 => x"8106bf38",
          9771 => x"82755f57",
          9772 => x"7652923d",
          9773 => x"f00551c1",
          9774 => x"f43f82b6",
          9775 => x"9808ff2e",
          9776 => x"d13882b6",
          9777 => x"9808812e",
          9778 => x"ce3882b6",
          9779 => x"98083070",
          9780 => x"82b69808",
          9781 => x"0780257a",
          9782 => x"0581197f",
          9783 => x"53595a54",
          9784 => x"98140877",
          9785 => x"26ca3880",
          9786 => x"f939a415",
          9787 => x"0882b698",
          9788 => x"08575875",
          9789 => x"98387752",
          9790 => x"81187d52",
          9791 => x"58ffbf8d",
          9792 => x"3f82b698",
          9793 => x"085b82b6",
          9794 => x"980880d6",
          9795 => x"387c7033",
          9796 => x"7712ff1a",
          9797 => x"5d525654",
          9798 => x"74822e09",
          9799 => x"81069e38",
          9800 => x"b41451ff",
          9801 => x"bbcb3f82",
          9802 => x"b6980883",
          9803 => x"ffff0670",
          9804 => x"30708025",
          9805 => x"1b821959",
          9806 => x"5b51549b",
          9807 => x"39b41451",
          9808 => x"ffbbc53f",
          9809 => x"82b69808",
          9810 => x"f00a0670",
          9811 => x"30708025",
          9812 => x"1b841959",
          9813 => x"5b515475",
          9814 => x"83ff067a",
          9815 => x"585679ff",
          9816 => x"9238787c",
          9817 => x"0c7c7990",
          9818 => x"120c8411",
          9819 => x"33810756",
          9820 => x"54748415",
          9821 => x"347a82b6",
          9822 => x"980c923d",
          9823 => x"0d04f93d",
          9824 => x"0d798a3d",
          9825 => x"fc055370",
          9826 => x"5257e3dd",
          9827 => x"3f82b698",
          9828 => x"085682b6",
          9829 => x"980881a8",
          9830 => x"38911733",
          9831 => x"567581a0",
          9832 => x"38901733",
          9833 => x"70812a70",
          9834 => x"81065155",
          9835 => x"55875573",
          9836 => x"802e818e",
          9837 => x"38941708",
          9838 => x"54738c18",
          9839 => x"08278180",
          9840 => x"38739b38",
          9841 => x"82b69808",
          9842 => x"53881708",
          9843 => x"527651c4",
          9844 => x"8c3f82b6",
          9845 => x"98087488",
          9846 => x"190c5680",
          9847 => x"c9399817",
          9848 => x"08527651",
          9849 => x"ffbfc63f",
          9850 => x"82b69808",
          9851 => x"ff2e0981",
          9852 => x"06833881",
          9853 => x"5682b698",
          9854 => x"08812e09",
          9855 => x"81068538",
          9856 => x"8256a339",
          9857 => x"75a03877",
          9858 => x"5482b698",
          9859 => x"08981508",
          9860 => x"27943898",
          9861 => x"17085382",
          9862 => x"b6980852",
          9863 => x"7651c3bd",
          9864 => x"3f82b698",
          9865 => x"08569417",
          9866 => x"088c180c",
          9867 => x"90173380",
          9868 => x"c0075473",
          9869 => x"90183475",
          9870 => x"802e8538",
          9871 => x"75911834",
          9872 => x"75557482",
          9873 => x"b6980c89",
          9874 => x"3d0d04e2",
          9875 => x"3d0d8253",
          9876 => x"a03dffa4",
          9877 => x"0552a13d",
          9878 => x"51dae43f",
          9879 => x"82b69808",
          9880 => x"5582b698",
          9881 => x"0881f538",
          9882 => x"7845a13d",
          9883 => x"0852953d",
          9884 => x"705258d1",
          9885 => x"ae3f82b6",
          9886 => x"98085582",
          9887 => x"b6980881",
          9888 => x"db380280",
          9889 => x"fb053370",
          9890 => x"852a7081",
          9891 => x"06515556",
          9892 => x"86557381",
          9893 => x"c7387598",
          9894 => x"2b548074",
          9895 => x"2481bd38",
          9896 => x"0280d605",
          9897 => x"33708106",
          9898 => x"58548755",
          9899 => x"7681ad38",
          9900 => x"6b527851",
          9901 => x"ccc53f82",
          9902 => x"b6980874",
          9903 => x"842a7081",
          9904 => x"06515556",
          9905 => x"73802e80",
          9906 => x"d4387854",
          9907 => x"82b69808",
          9908 => x"9415082e",
          9909 => x"81863873",
          9910 => x"5a82b698",
          9911 => x"085c7652",
          9912 => x"8a3d7052",
          9913 => x"54c7b53f",
          9914 => x"82b69808",
          9915 => x"5582b698",
          9916 => x"0880e938",
          9917 => x"82b69808",
          9918 => x"527351cc",
          9919 => x"e53f82b6",
          9920 => x"98085582",
          9921 => x"b6980886",
          9922 => x"38875580",
          9923 => x"cf3982b6",
          9924 => x"9808842e",
          9925 => x"883882b6",
          9926 => x"980880c0",
          9927 => x"387751ce",
          9928 => x"c23f82b6",
          9929 => x"980882b6",
          9930 => x"98083070",
          9931 => x"82b69808",
          9932 => x"07802551",
          9933 => x"55557580",
          9934 => x"2e943873",
          9935 => x"802e8f38",
          9936 => x"80537552",
          9937 => x"7751c195",
          9938 => x"3f82b698",
          9939 => x"0855748c",
          9940 => x"387851ff",
          9941 => x"bafe3f82",
          9942 => x"b6980855",
          9943 => x"7482b698",
          9944 => x"0ca03d0d",
          9945 => x"04e93d0d",
          9946 => x"8253993d",
          9947 => x"c005529a",
          9948 => x"3d51d8cb",
          9949 => x"3f82b698",
          9950 => x"085482b6",
          9951 => x"980882b0",
          9952 => x"38785e69",
          9953 => x"528e3d70",
          9954 => x"5258cf97",
          9955 => x"3f82b698",
          9956 => x"085482b6",
          9957 => x"98088638",
          9958 => x"88548294",
          9959 => x"3982b698",
          9960 => x"08842e09",
          9961 => x"81068288",
          9962 => x"380280df",
          9963 => x"05337085",
          9964 => x"2a810651",
          9965 => x"55865474",
          9966 => x"81f63878",
          9967 => x"5a74528a",
          9968 => x"3d705257",
          9969 => x"c1c33f82",
          9970 => x"b6980875",
          9971 => x"555682b6",
          9972 => x"98088338",
          9973 => x"875482b6",
          9974 => x"9808812e",
          9975 => x"09810683",
          9976 => x"38825482",
          9977 => x"b69808ff",
          9978 => x"2e098106",
          9979 => x"86388154",
          9980 => x"81b43973",
          9981 => x"81b03882",
          9982 => x"b6980852",
          9983 => x"7851c4a4",
          9984 => x"3f82b698",
          9985 => x"085482b6",
          9986 => x"9808819a",
          9987 => x"388b53a0",
          9988 => x"52b41951",
          9989 => x"ffb78c3f",
          9990 => x"7854ae0b",
          9991 => x"b4153478",
          9992 => x"54900bbf",
          9993 => x"15348288",
          9994 => x"b20a5280",
          9995 => x"ca1951ff",
          9996 => x"b69f3f75",
          9997 => x"5378b411",
          9998 => x"5351c9f8",
          9999 => x"3fa05378",
         10000 => x"b4115380",
         10001 => x"d40551ff",
         10002 => x"b6b63f78",
         10003 => x"54ae0b80",
         10004 => x"d515347f",
         10005 => x"537880d4",
         10006 => x"115351c9",
         10007 => x"d73f7854",
         10008 => x"810b8315",
         10009 => x"347751cb",
         10010 => x"a43f82b6",
         10011 => x"98085482",
         10012 => x"b69808b2",
         10013 => x"388288b2",
         10014 => x"0a526496",
         10015 => x"0551ffb5",
         10016 => x"d03f7553",
         10017 => x"64527851",
         10018 => x"c9aa3f64",
         10019 => x"54900b8b",
         10020 => x"15347854",
         10021 => x"810b8315",
         10022 => x"347851ff",
         10023 => x"b8b63f82",
         10024 => x"b6980854",
         10025 => x"8b398053",
         10026 => x"75527651",
         10027 => x"ffbeae3f",
         10028 => x"7382b698",
         10029 => x"0c993d0d",
         10030 => x"04da3d0d",
         10031 => x"a93d8405",
         10032 => x"51d2f13f",
         10033 => x"8253a83d",
         10034 => x"ff840552",
         10035 => x"a93d51d5",
         10036 => x"ee3f82b6",
         10037 => x"98085582",
         10038 => x"b6980882",
         10039 => x"d338784d",
         10040 => x"a93d0852",
         10041 => x"9d3d7052",
         10042 => x"58ccb83f",
         10043 => x"82b69808",
         10044 => x"5582b698",
         10045 => x"0882b938",
         10046 => x"02819b05",
         10047 => x"3381a006",
         10048 => x"54865573",
         10049 => x"82aa38a0",
         10050 => x"53a43d08",
         10051 => x"52a83dff",
         10052 => x"880551ff",
         10053 => x"b4ea3fac",
         10054 => x"53775292",
         10055 => x"3d705254",
         10056 => x"ffb4dd3f",
         10057 => x"aa3d0852",
         10058 => x"7351cbf7",
         10059 => x"3f82b698",
         10060 => x"085582b6",
         10061 => x"98089538",
         10062 => x"636f2e09",
         10063 => x"81068838",
         10064 => x"65a23d08",
         10065 => x"2e923888",
         10066 => x"5581e539",
         10067 => x"82b69808",
         10068 => x"842e0981",
         10069 => x"0681b838",
         10070 => x"7351c9b1",
         10071 => x"3f82b698",
         10072 => x"085582b6",
         10073 => x"980881c8",
         10074 => x"38685693",
         10075 => x"53a83dff",
         10076 => x"9505528d",
         10077 => x"1651ffb4",
         10078 => x"873f02af",
         10079 => x"05338b17",
         10080 => x"348b1633",
         10081 => x"70842a70",
         10082 => x"81065155",
         10083 => x"55738938",
         10084 => x"74a00754",
         10085 => x"738b1734",
         10086 => x"7854810b",
         10087 => x"8315348b",
         10088 => x"16337084",
         10089 => x"2a708106",
         10090 => x"51555573",
         10091 => x"802e80e5",
         10092 => x"386e642e",
         10093 => x"80df3875",
         10094 => x"527851c6",
         10095 => x"be3f82b6",
         10096 => x"98085278",
         10097 => x"51ffb7bb",
         10098 => x"3f825582",
         10099 => x"b6980880",
         10100 => x"2e80dd38",
         10101 => x"82b69808",
         10102 => x"527851ff",
         10103 => x"b5af3f82",
         10104 => x"b6980879",
         10105 => x"80d41158",
         10106 => x"585582b6",
         10107 => x"980880c0",
         10108 => x"38811633",
         10109 => x"5473ae2e",
         10110 => x"09810699",
         10111 => x"38635375",
         10112 => x"527651c6",
         10113 => x"af3f7854",
         10114 => x"810b8315",
         10115 => x"34873982",
         10116 => x"b698089c",
         10117 => x"387751c8",
         10118 => x"ca3f82b6",
         10119 => x"98085582",
         10120 => x"b698088c",
         10121 => x"387851ff",
         10122 => x"b5aa3f82",
         10123 => x"b6980855",
         10124 => x"7482b698",
         10125 => x"0ca83d0d",
         10126 => x"04ed3d0d",
         10127 => x"0280db05",
         10128 => x"33028405",
         10129 => x"80df0533",
         10130 => x"57578253",
         10131 => x"953dd005",
         10132 => x"52963d51",
         10133 => x"d2e93f82",
         10134 => x"b6980855",
         10135 => x"82b69808",
         10136 => x"80cf3878",
         10137 => x"5a655295",
         10138 => x"3dd40551",
         10139 => x"c9b53f82",
         10140 => x"b6980855",
         10141 => x"82b69808",
         10142 => x"b8380280",
         10143 => x"cf053381",
         10144 => x"a0065486",
         10145 => x"5573aa38",
         10146 => x"75a70661",
         10147 => x"71098b12",
         10148 => x"3371067a",
         10149 => x"74060751",
         10150 => x"57555674",
         10151 => x"8b153478",
         10152 => x"54810b83",
         10153 => x"15347851",
         10154 => x"ffb4a93f",
         10155 => x"82b69808",
         10156 => x"557482b6",
         10157 => x"980c953d",
         10158 => x"0d04ef3d",
         10159 => x"0d645682",
         10160 => x"53933dd0",
         10161 => x"0552943d",
         10162 => x"51d1f43f",
         10163 => x"82b69808",
         10164 => x"5582b698",
         10165 => x"0880cb38",
         10166 => x"76586352",
         10167 => x"933dd405",
         10168 => x"51c8c03f",
         10169 => x"82b69808",
         10170 => x"5582b698",
         10171 => x"08b43802",
         10172 => x"80c70533",
         10173 => x"81a00654",
         10174 => x"865573a6",
         10175 => x"38841622",
         10176 => x"86172271",
         10177 => x"902b0753",
         10178 => x"54961f51",
         10179 => x"ffb0c23f",
         10180 => x"7654810b",
         10181 => x"83153476",
         10182 => x"51ffb3b8",
         10183 => x"3f82b698",
         10184 => x"08557482",
         10185 => x"b6980c93",
         10186 => x"3d0d04ea",
         10187 => x"3d0d696b",
         10188 => x"5c5a8053",
         10189 => x"983dd005",
         10190 => x"52993d51",
         10191 => x"d1813f82",
         10192 => x"b6980882",
         10193 => x"b6980830",
         10194 => x"7082b698",
         10195 => x"08078025",
         10196 => x"51555779",
         10197 => x"802e8185",
         10198 => x"38817075",
         10199 => x"06555573",
         10200 => x"802e80f9",
         10201 => x"387b5d80",
         10202 => x"5f80528d",
         10203 => x"3d705254",
         10204 => x"ffbea93f",
         10205 => x"82b69808",
         10206 => x"5782b698",
         10207 => x"0880d138",
         10208 => x"74527351",
         10209 => x"c3dc3f82",
         10210 => x"b6980857",
         10211 => x"82b69808",
         10212 => x"bf3882b6",
         10213 => x"980882b6",
         10214 => x"9808655b",
         10215 => x"59567818",
         10216 => x"81197b18",
         10217 => x"56595574",
         10218 => x"33743481",
         10219 => x"16568a78",
         10220 => x"27ec388b",
         10221 => x"56751a54",
         10222 => x"80743475",
         10223 => x"802e9e38",
         10224 => x"ff16701b",
         10225 => x"70335155",
         10226 => x"5673a02e",
         10227 => x"e8388e39",
         10228 => x"76842e09",
         10229 => x"81068638",
         10230 => x"807a3480",
         10231 => x"57763070",
         10232 => x"78078025",
         10233 => x"51547a80",
         10234 => x"2e80c138",
         10235 => x"73802ebc",
         10236 => x"387ba011",
         10237 => x"085351ff",
         10238 => x"b1933f82",
         10239 => x"b6980857",
         10240 => x"82b69808",
         10241 => x"a7387b70",
         10242 => x"33555580",
         10243 => x"c3567383",
         10244 => x"2e8b3880",
         10245 => x"e4567384",
         10246 => x"2e8338a7",
         10247 => x"567515b4",
         10248 => x"0551ffad",
         10249 => x"e33f82b6",
         10250 => x"98087b0c",
         10251 => x"7682b698",
         10252 => x"0c983d0d",
         10253 => x"04e63d0d",
         10254 => x"82539c3d",
         10255 => x"ffb80552",
         10256 => x"9d3d51ce",
         10257 => x"fa3f82b6",
         10258 => x"980882b6",
         10259 => x"98085654",
         10260 => x"82b69808",
         10261 => x"8398388b",
         10262 => x"53a0528b",
         10263 => x"3d705259",
         10264 => x"ffaec03f",
         10265 => x"736d7033",
         10266 => x"7081ff06",
         10267 => x"52575557",
         10268 => x"9f742781",
         10269 => x"bc387858",
         10270 => x"7481ff06",
         10271 => x"6d81054e",
         10272 => x"705255ff",
         10273 => x"af893f82",
         10274 => x"b6980880",
         10275 => x"2ea5386c",
         10276 => x"70337053",
         10277 => x"5754ffae",
         10278 => x"fd3f82b6",
         10279 => x"9808802e",
         10280 => x"8d387488",
         10281 => x"2b76076d",
         10282 => x"81054e55",
         10283 => x"863982b6",
         10284 => x"980855ff",
         10285 => x"9f157083",
         10286 => x"ffff0651",
         10287 => x"54739926",
         10288 => x"8a38e015",
         10289 => x"7083ffff",
         10290 => x"06565480",
         10291 => x"ff752787",
         10292 => x"3882aee0",
         10293 => x"15335574",
         10294 => x"802ea338",
         10295 => x"745282b0",
         10296 => x"e051ffae",
         10297 => x"893f82b6",
         10298 => x"98089338",
         10299 => x"81ff7527",
         10300 => x"88387689",
         10301 => x"2688388b",
         10302 => x"398a7727",
         10303 => x"86388655",
         10304 => x"81ec3981",
         10305 => x"ff75278f",
         10306 => x"3874882a",
         10307 => x"54737870",
         10308 => x"81055a34",
         10309 => x"81175774",
         10310 => x"78708105",
         10311 => x"5a348117",
         10312 => x"6d703370",
         10313 => x"81ff0652",
         10314 => x"57555773",
         10315 => x"9f26fec8",
         10316 => x"388b3d33",
         10317 => x"54865573",
         10318 => x"81e52e81",
         10319 => x"b1387680",
         10320 => x"2e993802",
         10321 => x"a7055576",
         10322 => x"15703351",
         10323 => x"5473a02e",
         10324 => x"09810687",
         10325 => x"38ff1757",
         10326 => x"76ed3879",
         10327 => x"41804380",
         10328 => x"52913d70",
         10329 => x"5255ffba",
         10330 => x"b33f82b6",
         10331 => x"98085482",
         10332 => x"b6980880",
         10333 => x"f7388152",
         10334 => x"7451ffbf",
         10335 => x"e53f82b6",
         10336 => x"98085482",
         10337 => x"b698088d",
         10338 => x"387680c4",
         10339 => x"386754e5",
         10340 => x"743480c6",
         10341 => x"3982b698",
         10342 => x"08842e09",
         10343 => x"810680cc",
         10344 => x"38805476",
         10345 => x"742e80c4",
         10346 => x"38815274",
         10347 => x"51ffbdb0",
         10348 => x"3f82b698",
         10349 => x"085482b6",
         10350 => x"9808b138",
         10351 => x"a05382b6",
         10352 => x"98085267",
         10353 => x"51ffabdb",
         10354 => x"3f675488",
         10355 => x"0b8b1534",
         10356 => x"8b537852",
         10357 => x"6751ffab",
         10358 => x"a73f7954",
         10359 => x"810b8315",
         10360 => x"347951ff",
         10361 => x"adee3f82",
         10362 => x"b6980854",
         10363 => x"73557482",
         10364 => x"b6980c9c",
         10365 => x"3d0d04f2",
         10366 => x"3d0d6062",
         10367 => x"02880580",
         10368 => x"cb053393",
         10369 => x"3dfc0555",
         10370 => x"7254405e",
         10371 => x"5ad2da3f",
         10372 => x"82b69808",
         10373 => x"5882b698",
         10374 => x"0882bd38",
         10375 => x"911a3358",
         10376 => x"7782b538",
         10377 => x"7c802e97",
         10378 => x"388c1a08",
         10379 => x"59789038",
         10380 => x"901a3370",
         10381 => x"812a7081",
         10382 => x"06515555",
         10383 => x"73903887",
         10384 => x"54829739",
         10385 => x"82588290",
         10386 => x"39815882",
         10387 => x"8b397e8a",
         10388 => x"11227089",
         10389 => x"2b70557f",
         10390 => x"54565656",
         10391 => x"fec2a43f",
         10392 => x"ff147d06",
         10393 => x"70307072",
         10394 => x"079f2a82",
         10395 => x"b6980805",
         10396 => x"8c19087c",
         10397 => x"405a5d55",
         10398 => x"55817727",
         10399 => x"88389816",
         10400 => x"08772683",
         10401 => x"38825776",
         10402 => x"77565980",
         10403 => x"56745279",
         10404 => x"51ffae99",
         10405 => x"3f81157f",
         10406 => x"55559814",
         10407 => x"08752683",
         10408 => x"38825582",
         10409 => x"b6980881",
         10410 => x"2eff9938",
         10411 => x"82b69808",
         10412 => x"ff2eff95",
         10413 => x"3882b698",
         10414 => x"088e3881",
         10415 => x"1656757b",
         10416 => x"2e098106",
         10417 => x"87389339",
         10418 => x"74598056",
         10419 => x"74772e09",
         10420 => x"8106ffb9",
         10421 => x"38875880",
         10422 => x"ff397d80",
         10423 => x"2eba3878",
         10424 => x"7b55557a",
         10425 => x"802eb438",
         10426 => x"81155673",
         10427 => x"812e0981",
         10428 => x"068338ff",
         10429 => x"56755374",
         10430 => x"527e51ff",
         10431 => x"afa83f82",
         10432 => x"b6980858",
         10433 => x"82b69808",
         10434 => x"80ce3874",
         10435 => x"8116ff16",
         10436 => x"56565c73",
         10437 => x"d3388439",
         10438 => x"ff195c7e",
         10439 => x"7c8c120c",
         10440 => x"557d802e",
         10441 => x"b3387888",
         10442 => x"1b0c7c8c",
         10443 => x"1b0c901a",
         10444 => x"3380c007",
         10445 => x"5473901b",
         10446 => x"34981508",
         10447 => x"fe059016",
         10448 => x"08575475",
         10449 => x"74269138",
         10450 => x"757b3190",
         10451 => x"160c8415",
         10452 => x"33810754",
         10453 => x"73841634",
         10454 => x"77547382",
         10455 => x"b6980c90",
         10456 => x"3d0d04e9",
         10457 => x"3d0d6b6d",
         10458 => x"02880580",
         10459 => x"eb05339d",
         10460 => x"3d545a5c",
         10461 => x"59c5bd3f",
         10462 => x"8b56800b",
         10463 => x"82b69808",
         10464 => x"248bf838",
         10465 => x"82b69808",
         10466 => x"842982cd",
         10467 => x"d0057008",
         10468 => x"51557480",
         10469 => x"2e843880",
         10470 => x"753482b6",
         10471 => x"980881ff",
         10472 => x"065f8152",
         10473 => x"7e51ffa0",
         10474 => x"d03f82b6",
         10475 => x"980881ff",
         10476 => x"06708106",
         10477 => x"56578356",
         10478 => x"748bc038",
         10479 => x"76822a70",
         10480 => x"81065155",
         10481 => x"8a56748b",
         10482 => x"b238993d",
         10483 => x"fc055383",
         10484 => x"527e51ff",
         10485 => x"a4f03f82",
         10486 => x"b6980899",
         10487 => x"38675574",
         10488 => x"802e9238",
         10489 => x"74828080",
         10490 => x"268b38ff",
         10491 => x"15750655",
         10492 => x"74802e83",
         10493 => x"38814878",
         10494 => x"802e8738",
         10495 => x"84807926",
         10496 => x"92387881",
         10497 => x"800a268b",
         10498 => x"38ff1979",
         10499 => x"06557480",
         10500 => x"2e863893",
         10501 => x"568ae439",
         10502 => x"78892a6e",
         10503 => x"892a7089",
         10504 => x"2b775948",
         10505 => x"43597a83",
         10506 => x"38815661",
         10507 => x"30708025",
         10508 => x"77075155",
         10509 => x"9156748a",
         10510 => x"c238993d",
         10511 => x"f8055381",
         10512 => x"527e51ff",
         10513 => x"a4803f81",
         10514 => x"5682b698",
         10515 => x"088aac38",
         10516 => x"77832a70",
         10517 => x"770682b6",
         10518 => x"98084356",
         10519 => x"45748338",
         10520 => x"bf416655",
         10521 => x"8e566075",
         10522 => x"268a9038",
         10523 => x"74613170",
         10524 => x"485580ff",
         10525 => x"75278a83",
         10526 => x"38935678",
         10527 => x"81802689",
         10528 => x"fa387781",
         10529 => x"2a708106",
         10530 => x"56437480",
         10531 => x"2e953877",
         10532 => x"87065574",
         10533 => x"822e838d",
         10534 => x"38778106",
         10535 => x"5574802e",
         10536 => x"83833877",
         10537 => x"81065593",
         10538 => x"56825e74",
         10539 => x"802e89cb",
         10540 => x"38785a7d",
         10541 => x"832e0981",
         10542 => x"0680e138",
         10543 => x"78ae3866",
         10544 => x"912a5781",
         10545 => x"0b82b184",
         10546 => x"22565a74",
         10547 => x"802e9d38",
         10548 => x"74772698",
         10549 => x"3882b184",
         10550 => x"56791082",
         10551 => x"17702257",
         10552 => x"575a7480",
         10553 => x"2e863876",
         10554 => x"7527ee38",
         10555 => x"79526651",
         10556 => x"febd903f",
         10557 => x"82b69808",
         10558 => x"84298487",
         10559 => x"0570892a",
         10560 => x"5e55a05c",
         10561 => x"800b82b6",
         10562 => x"9808fc80",
         10563 => x"8a055644",
         10564 => x"fdfff00a",
         10565 => x"752780ec",
         10566 => x"3888d339",
         10567 => x"78ae3866",
         10568 => x"8c2a5781",
         10569 => x"0b82b0f4",
         10570 => x"22565a74",
         10571 => x"802e9d38",
         10572 => x"74772698",
         10573 => x"3882b0f4",
         10574 => x"56791082",
         10575 => x"17702257",
         10576 => x"575a7480",
         10577 => x"2e863876",
         10578 => x"7527ee38",
         10579 => x"79526651",
         10580 => x"febcb03f",
         10581 => x"82b69808",
         10582 => x"10840557",
         10583 => x"82b69808",
         10584 => x"9ff52696",
         10585 => x"38810b82",
         10586 => x"b6980810",
         10587 => x"82b69808",
         10588 => x"05711172",
         10589 => x"2a830559",
         10590 => x"565e83ff",
         10591 => x"17892a5d",
         10592 => x"815ca044",
         10593 => x"601c7d11",
         10594 => x"65056970",
         10595 => x"12ff0571",
         10596 => x"30707206",
         10597 => x"74315c52",
         10598 => x"59575940",
         10599 => x"7d832e09",
         10600 => x"81068938",
         10601 => x"761c6018",
         10602 => x"415c8439",
         10603 => x"761d5d79",
         10604 => x"90291870",
         10605 => x"62316858",
         10606 => x"51557476",
         10607 => x"2687af38",
         10608 => x"757c317d",
         10609 => x"317a5370",
         10610 => x"65315255",
         10611 => x"febbb43f",
         10612 => x"82b69808",
         10613 => x"587d832e",
         10614 => x"0981069b",
         10615 => x"3882b698",
         10616 => x"0883fff5",
         10617 => x"2680dd38",
         10618 => x"78878338",
         10619 => x"79812a59",
         10620 => x"78fdbe38",
         10621 => x"86f8397d",
         10622 => x"822e0981",
         10623 => x"0680c538",
         10624 => x"83fff50b",
         10625 => x"82b69808",
         10626 => x"27a03878",
         10627 => x"8f38791a",
         10628 => x"557480c0",
         10629 => x"26863874",
         10630 => x"59fd9639",
         10631 => x"62810655",
         10632 => x"74802e8f",
         10633 => x"38835efd",
         10634 => x"883982b6",
         10635 => x"98089ff5",
         10636 => x"26923878",
         10637 => x"86b83879",
         10638 => x"1a598180",
         10639 => x"7927fcf1",
         10640 => x"3886ab39",
         10641 => x"80557d81",
         10642 => x"2e098106",
         10643 => x"83387d55",
         10644 => x"9ff57827",
         10645 => x"8b387481",
         10646 => x"06558e56",
         10647 => x"74869c38",
         10648 => x"84805380",
         10649 => x"527a51ff",
         10650 => x"a2b93f8b",
         10651 => x"5382af9c",
         10652 => x"527a51ff",
         10653 => x"a28a3f84",
         10654 => x"80528b1b",
         10655 => x"51ffa1b3",
         10656 => x"3f798d1c",
         10657 => x"347b83ff",
         10658 => x"ff06528e",
         10659 => x"1b51ffa1",
         10660 => x"a23f810b",
         10661 => x"901c347d",
         10662 => x"83327030",
         10663 => x"70962a84",
         10664 => x"80065451",
         10665 => x"55911b51",
         10666 => x"ffa1883f",
         10667 => x"66557483",
         10668 => x"ffff2690",
         10669 => x"387483ff",
         10670 => x"ff065293",
         10671 => x"1b51ffa0",
         10672 => x"f23f8a39",
         10673 => x"7452a01b",
         10674 => x"51ffa185",
         10675 => x"3ff80b95",
         10676 => x"1c34bf52",
         10677 => x"981b51ff",
         10678 => x"a0d93f81",
         10679 => x"ff529a1b",
         10680 => x"51ffa0cf",
         10681 => x"3f60529c",
         10682 => x"1b51ffa0",
         10683 => x"e43f7d83",
         10684 => x"2e098106",
         10685 => x"80cb3882",
         10686 => x"88b20a52",
         10687 => x"80c31b51",
         10688 => x"ffa0ce3f",
         10689 => x"7c52a41b",
         10690 => x"51ffa0c5",
         10691 => x"3f8252ac",
         10692 => x"1b51ffa0",
         10693 => x"bc3f8152",
         10694 => x"b01b51ff",
         10695 => x"a0953f86",
         10696 => x"52b21b51",
         10697 => x"ffa08c3f",
         10698 => x"ff800b80",
         10699 => x"c01c34a9",
         10700 => x"0b80c21c",
         10701 => x"34935382",
         10702 => x"afa85280",
         10703 => x"c71b51ae",
         10704 => x"398288b2",
         10705 => x"0a52a71b",
         10706 => x"51ffa085",
         10707 => x"3f7c83ff",
         10708 => x"ff065296",
         10709 => x"1b51ff9f",
         10710 => x"da3fff80",
         10711 => x"0ba41c34",
         10712 => x"a90ba61c",
         10713 => x"34935382",
         10714 => x"afbc52ab",
         10715 => x"1b51ffa0",
         10716 => x"8f3f82d4",
         10717 => x"d55283fe",
         10718 => x"1b705259",
         10719 => x"ff9fb43f",
         10720 => x"81546053",
         10721 => x"7a527e51",
         10722 => x"ff9bd73f",
         10723 => x"815682b6",
         10724 => x"980883e7",
         10725 => x"387d832e",
         10726 => x"09810680",
         10727 => x"ee387554",
         10728 => x"60860553",
         10729 => x"7a527e51",
         10730 => x"ff9bb73f",
         10731 => x"84805380",
         10732 => x"527a51ff",
         10733 => x"9fed3f84",
         10734 => x"8b85a4d2",
         10735 => x"527a51ff",
         10736 => x"9f8f3f86",
         10737 => x"8a85e4f2",
         10738 => x"5283e41b",
         10739 => x"51ff9f81",
         10740 => x"3fff1852",
         10741 => x"83e81b51",
         10742 => x"ff9ef63f",
         10743 => x"825283ec",
         10744 => x"1b51ff9e",
         10745 => x"ec3f82d4",
         10746 => x"d5527851",
         10747 => x"ff9ec43f",
         10748 => x"75546087",
         10749 => x"05537a52",
         10750 => x"7e51ff9a",
         10751 => x"e53f7554",
         10752 => x"6016537a",
         10753 => x"527e51ff",
         10754 => x"9ad83f65",
         10755 => x"5380527a",
         10756 => x"51ff9f8f",
         10757 => x"3f7f5680",
         10758 => x"587d832e",
         10759 => x"0981069a",
         10760 => x"38f8527a",
         10761 => x"51ff9ea9",
         10762 => x"3fff5284",
         10763 => x"1b51ff9e",
         10764 => x"a03ff00a",
         10765 => x"52881b51",
         10766 => x"913987ff",
         10767 => x"fff8557d",
         10768 => x"812e8338",
         10769 => x"f8557452",
         10770 => x"7a51ff9e",
         10771 => x"843f7c55",
         10772 => x"61577462",
         10773 => x"26833874",
         10774 => x"57765475",
         10775 => x"537a527e",
         10776 => x"51ff99fe",
         10777 => x"3f82b698",
         10778 => x"08828738",
         10779 => x"84805382",
         10780 => x"b6980852",
         10781 => x"7a51ff9e",
         10782 => x"aa3f7616",
         10783 => x"75783156",
         10784 => x"5674cd38",
         10785 => x"81185877",
         10786 => x"802eff8d",
         10787 => x"3879557d",
         10788 => x"832e8338",
         10789 => x"63556157",
         10790 => x"74622683",
         10791 => x"38745776",
         10792 => x"5475537a",
         10793 => x"527e51ff",
         10794 => x"99b83f82",
         10795 => x"b6980881",
         10796 => x"c1387616",
         10797 => x"75783156",
         10798 => x"5674db38",
         10799 => x"8c567d83",
         10800 => x"2e933886",
         10801 => x"566683ff",
         10802 => x"ff268a38",
         10803 => x"84567d82",
         10804 => x"2e833881",
         10805 => x"56648106",
         10806 => x"587780fe",
         10807 => x"38848053",
         10808 => x"77527a51",
         10809 => x"ff9dbc3f",
         10810 => x"82d4d552",
         10811 => x"7851ff9c",
         10812 => x"c23f83be",
         10813 => x"1b557775",
         10814 => x"34810b81",
         10815 => x"1634810b",
         10816 => x"82163477",
         10817 => x"83163475",
         10818 => x"84163460",
         10819 => x"67055680",
         10820 => x"fdc15275",
         10821 => x"51feb4eb",
         10822 => x"3ffe0b85",
         10823 => x"163482b6",
         10824 => x"9808822a",
         10825 => x"bf075675",
         10826 => x"86163482",
         10827 => x"b6980887",
         10828 => x"16346052",
         10829 => x"83c61b51",
         10830 => x"ff9c963f",
         10831 => x"665283ca",
         10832 => x"1b51ff9c",
         10833 => x"8c3f8154",
         10834 => x"77537a52",
         10835 => x"7e51ff98",
         10836 => x"913f8156",
         10837 => x"82b69808",
         10838 => x"a2388053",
         10839 => x"80527e51",
         10840 => x"ff99e33f",
         10841 => x"815682b6",
         10842 => x"98089038",
         10843 => x"89398e56",
         10844 => x"8a398156",
         10845 => x"863982b6",
         10846 => x"98085675",
         10847 => x"82b6980c",
         10848 => x"993d0d04",
         10849 => x"f53d0d7d",
         10850 => x"605b5980",
         10851 => x"7960ff05",
         10852 => x"5a575776",
         10853 => x"7825b438",
         10854 => x"8d3df811",
         10855 => x"55558153",
         10856 => x"fc155279",
         10857 => x"51c9dc3f",
         10858 => x"7a812e09",
         10859 => x"81069c38",
         10860 => x"8c3d3355",
         10861 => x"748d2edb",
         10862 => x"38747670",
         10863 => x"81055834",
         10864 => x"81175774",
         10865 => x"8a2e0981",
         10866 => x"06c93880",
         10867 => x"76347855",
         10868 => x"76833876",
         10869 => x"557482b6",
         10870 => x"980c8d3d",
         10871 => x"0d04f73d",
         10872 => x"0d7b0284",
         10873 => x"05b30533",
         10874 => x"5957778a",
         10875 => x"2e098106",
         10876 => x"87388d52",
         10877 => x"7651e73f",
         10878 => x"84170856",
         10879 => x"807624be",
         10880 => x"38881708",
         10881 => x"77178c05",
         10882 => x"56597775",
         10883 => x"34811656",
         10884 => x"bb7625a1",
         10885 => x"388b3dfc",
         10886 => x"05547553",
         10887 => x"8c175276",
         10888 => x"0851cbdc",
         10889 => x"3f797632",
         10890 => x"70307072",
         10891 => x"079f2a70",
         10892 => x"30535156",
         10893 => x"56758418",
         10894 => x"0c811988",
         10895 => x"180c8b3d",
         10896 => x"0d04f93d",
         10897 => x"0d798411",
         10898 => x"08565680",
         10899 => x"7524a738",
         10900 => x"893dfc05",
         10901 => x"5474538c",
         10902 => x"16527508",
         10903 => x"51cba13f",
         10904 => x"82b69808",
         10905 => x"91388416",
         10906 => x"08782e09",
         10907 => x"81068738",
         10908 => x"88160855",
         10909 => x"8339ff55",
         10910 => x"7482b698",
         10911 => x"0c893d0d",
         10912 => x"04fd3d0d",
         10913 => x"755480cc",
         10914 => x"53805273",
         10915 => x"51ff9a93",
         10916 => x"3f76740c",
         10917 => x"853d0d04",
         10918 => x"ea3d0d02",
         10919 => x"80e30533",
         10920 => x"6a53863d",
         10921 => x"70535454",
         10922 => x"d83f7352",
         10923 => x"7251feae",
         10924 => x"3f7251ff",
         10925 => x"8d3f983d",
         10926 => x"0d040000",
         10927 => x"00ffffff",
         10928 => x"ff00ffff",
         10929 => x"ffff00ff",
         10930 => x"ffffff00",
         10931 => x"00002baa",
         10932 => x"00002b2e",
         10933 => x"00002b35",
         10934 => x"00002b3c",
         10935 => x"00002b43",
         10936 => x"00002b4a",
         10937 => x"00002b51",
         10938 => x"00002b58",
         10939 => x"00002b5f",
         10940 => x"00002b66",
         10941 => x"00002b6d",
         10942 => x"00002b74",
         10943 => x"00002b7a",
         10944 => x"00002b80",
         10945 => x"00002b86",
         10946 => x"00002b8c",
         10947 => x"00002b92",
         10948 => x"00002b98",
         10949 => x"00002b9e",
         10950 => x"00002ba4",
         10951 => x"00004171",
         10952 => x"00004177",
         10953 => x"0000417d",
         10954 => x"00004183",
         10955 => x"00004189",
         10956 => x"00004767",
         10957 => x"00004867",
         10958 => x"00004978",
         10959 => x"00004bd0",
         10960 => x"0000484f",
         10961 => x"0000463c",
         10962 => x"00004a40",
         10963 => x"00004ba1",
         10964 => x"00004a83",
         10965 => x"00004b19",
         10966 => x"00004a9f",
         10967 => x"00004922",
         10968 => x"0000463c",
         10969 => x"00004978",
         10970 => x"000049a1",
         10971 => x"00004a40",
         10972 => x"0000463c",
         10973 => x"0000463c",
         10974 => x"00004a9f",
         10975 => x"00004b19",
         10976 => x"00004ba1",
         10977 => x"00004bd0",
         10978 => x"00000e31",
         10979 => x"0000171a",
         10980 => x"0000171a",
         10981 => x"00000e60",
         10982 => x"0000171a",
         10983 => x"0000171a",
         10984 => x"0000171a",
         10985 => x"0000171a",
         10986 => x"0000171a",
         10987 => x"0000171a",
         10988 => x"0000171a",
         10989 => x"00000e1d",
         10990 => x"0000171a",
         10991 => x"00000e48",
         10992 => x"00000e78",
         10993 => x"0000171a",
         10994 => x"0000171a",
         10995 => x"0000171a",
         10996 => x"0000171a",
         10997 => x"0000171a",
         10998 => x"0000171a",
         10999 => x"0000171a",
         11000 => x"0000171a",
         11001 => x"0000171a",
         11002 => x"0000171a",
         11003 => x"0000171a",
         11004 => x"0000171a",
         11005 => x"0000171a",
         11006 => x"0000171a",
         11007 => x"0000171a",
         11008 => x"0000171a",
         11009 => x"0000171a",
         11010 => x"0000171a",
         11011 => x"0000171a",
         11012 => x"0000171a",
         11013 => x"0000171a",
         11014 => x"0000171a",
         11015 => x"0000171a",
         11016 => x"0000171a",
         11017 => x"0000171a",
         11018 => x"0000171a",
         11019 => x"0000171a",
         11020 => x"0000171a",
         11021 => x"0000171a",
         11022 => x"0000171a",
         11023 => x"0000171a",
         11024 => x"0000171a",
         11025 => x"0000171a",
         11026 => x"0000171a",
         11027 => x"0000171a",
         11028 => x"0000171a",
         11029 => x"00000fa8",
         11030 => x"0000171a",
         11031 => x"0000171a",
         11032 => x"0000171a",
         11033 => x"0000171a",
         11034 => x"00001116",
         11035 => x"0000171a",
         11036 => x"0000171a",
         11037 => x"0000171a",
         11038 => x"0000171a",
         11039 => x"0000171a",
         11040 => x"0000171a",
         11041 => x"0000171a",
         11042 => x"0000171a",
         11043 => x"0000171a",
         11044 => x"0000171a",
         11045 => x"00000ed8",
         11046 => x"0000103f",
         11047 => x"00000eaf",
         11048 => x"00000eaf",
         11049 => x"00000eaf",
         11050 => x"0000171a",
         11051 => x"0000103f",
         11052 => x"0000171a",
         11053 => x"0000171a",
         11054 => x"00000e98",
         11055 => x"0000171a",
         11056 => x"0000171a",
         11057 => x"000010ec",
         11058 => x"000010f7",
         11059 => x"0000171a",
         11060 => x"0000171a",
         11061 => x"00000f11",
         11062 => x"0000171a",
         11063 => x"0000111f",
         11064 => x"0000171a",
         11065 => x"0000171a",
         11066 => x"00001116",
         11067 => x"64696e69",
         11068 => x"74000000",
         11069 => x"64696f63",
         11070 => x"746c0000",
         11071 => x"66696e69",
         11072 => x"74000000",
         11073 => x"666c6f61",
         11074 => x"64000000",
         11075 => x"66657865",
         11076 => x"63000000",
         11077 => x"6d636c65",
         11078 => x"61720000",
         11079 => x"6d636f70",
         11080 => x"79000000",
         11081 => x"6d646966",
         11082 => x"66000000",
         11083 => x"6d64756d",
         11084 => x"70000000",
         11085 => x"6d656200",
         11086 => x"6d656800",
         11087 => x"6d657700",
         11088 => x"68696400",
         11089 => x"68696500",
         11090 => x"68666400",
         11091 => x"68666500",
         11092 => x"63616c6c",
         11093 => x"00000000",
         11094 => x"6a6d7000",
         11095 => x"72657374",
         11096 => x"61727400",
         11097 => x"72657365",
         11098 => x"74000000",
         11099 => x"696e666f",
         11100 => x"00000000",
         11101 => x"74657374",
         11102 => x"00000000",
         11103 => x"74626173",
         11104 => x"69630000",
         11105 => x"6d626173",
         11106 => x"69630000",
         11107 => x"6b696c6f",
         11108 => x"00000000",
         11109 => x"65640000",
         11110 => x"4469736b",
         11111 => x"20457272",
         11112 => x"6f720000",
         11113 => x"496e7465",
         11114 => x"726e616c",
         11115 => x"20657272",
         11116 => x"6f722e00",
         11117 => x"4469736b",
         11118 => x"206e6f74",
         11119 => x"20726561",
         11120 => x"64792e00",
         11121 => x"4e6f2066",
         11122 => x"696c6520",
         11123 => x"666f756e",
         11124 => x"642e0000",
         11125 => x"4e6f2070",
         11126 => x"61746820",
         11127 => x"666f756e",
         11128 => x"642e0000",
         11129 => x"496e7661",
         11130 => x"6c696420",
         11131 => x"66696c65",
         11132 => x"6e616d65",
         11133 => x"2e000000",
         11134 => x"41636365",
         11135 => x"73732064",
         11136 => x"656e6965",
         11137 => x"642e0000",
         11138 => x"46696c65",
         11139 => x"20616c72",
         11140 => x"65616479",
         11141 => x"20657869",
         11142 => x"7374732e",
         11143 => x"00000000",
         11144 => x"46696c65",
         11145 => x"2068616e",
         11146 => x"646c6520",
         11147 => x"696e7661",
         11148 => x"6c69642e",
         11149 => x"00000000",
         11150 => x"53442069",
         11151 => x"73207772",
         11152 => x"69746520",
         11153 => x"70726f74",
         11154 => x"65637465",
         11155 => x"642e0000",
         11156 => x"44726976",
         11157 => x"65206e75",
         11158 => x"6d626572",
         11159 => x"20697320",
         11160 => x"696e7661",
         11161 => x"6c69642e",
         11162 => x"00000000",
         11163 => x"4469736b",
         11164 => x"206e6f74",
         11165 => x"20656e61",
         11166 => x"626c6564",
         11167 => x"2e000000",
         11168 => x"4e6f2063",
         11169 => x"6f6d7061",
         11170 => x"7469626c",
         11171 => x"65206669",
         11172 => x"6c657379",
         11173 => x"7374656d",
         11174 => x"20666f75",
         11175 => x"6e64206f",
         11176 => x"6e206469",
         11177 => x"736b2e00",
         11178 => x"466f726d",
         11179 => x"61742061",
         11180 => x"626f7274",
         11181 => x"65642e00",
         11182 => x"54696d65",
         11183 => x"6f75742c",
         11184 => x"206f7065",
         11185 => x"72617469",
         11186 => x"6f6e2063",
         11187 => x"616e6365",
         11188 => x"6c6c6564",
         11189 => x"2e000000",
         11190 => x"46696c65",
         11191 => x"20697320",
         11192 => x"6c6f636b",
         11193 => x"65642e00",
         11194 => x"496e7375",
         11195 => x"66666963",
         11196 => x"69656e74",
         11197 => x"206d656d",
         11198 => x"6f72792e",
         11199 => x"00000000",
         11200 => x"546f6f20",
         11201 => x"6d616e79",
         11202 => x"206f7065",
         11203 => x"6e206669",
         11204 => x"6c65732e",
         11205 => x"00000000",
         11206 => x"50617261",
         11207 => x"6d657465",
         11208 => x"72732069",
         11209 => x"6e636f72",
         11210 => x"72656374",
         11211 => x"2e000000",
         11212 => x"53756363",
         11213 => x"6573732e",
         11214 => x"00000000",
         11215 => x"556e6b6e",
         11216 => x"6f776e20",
         11217 => x"6572726f",
         11218 => x"722e0000",
         11219 => x"0a256c75",
         11220 => x"20627974",
         11221 => x"65732025",
         11222 => x"73206174",
         11223 => x"20256c75",
         11224 => x"20627974",
         11225 => x"65732f73",
         11226 => x"65632e0a",
         11227 => x"00000000",
         11228 => x"72656164",
         11229 => x"00000000",
         11230 => x"303d2530",
         11231 => x"386c782c",
         11232 => x"20313d25",
         11233 => x"30386c78",
         11234 => x"2c20323d",
         11235 => x"2530386c",
         11236 => x"782c205f",
         11237 => x"494f423d",
         11238 => x"2530386c",
         11239 => x"78202530",
         11240 => x"386c7820",
         11241 => x"2530386c",
         11242 => x"780a0000",
         11243 => x"2530386c",
         11244 => x"58000000",
         11245 => x"3a202000",
         11246 => x"25303458",
         11247 => x"00000000",
         11248 => x"20202020",
         11249 => x"20202020",
         11250 => x"00000000",
         11251 => x"25303258",
         11252 => x"00000000",
         11253 => x"20200000",
         11254 => x"207c0000",
         11255 => x"7c000000",
         11256 => x"7a4f5300",
         11257 => x"0a2a2a20",
         11258 => x"25732028",
         11259 => x"00000000",
         11260 => x"30322f30",
         11261 => x"352f3230",
         11262 => x"32300000",
         11263 => x"76312e30",
         11264 => x"32000000",
         11265 => x"205a5055",
         11266 => x"2c207265",
         11267 => x"76202530",
         11268 => x"32782920",
         11269 => x"25732025",
         11270 => x"73202a2a",
         11271 => x"0a0a0000",
         11272 => x"5a505520",
         11273 => x"496e7465",
         11274 => x"72727570",
         11275 => x"74204861",
         11276 => x"6e646c65",
         11277 => x"72000000",
         11278 => x"54696d65",
         11279 => x"7220696e",
         11280 => x"74657272",
         11281 => x"75707400",
         11282 => x"50533220",
         11283 => x"696e7465",
         11284 => x"72727570",
         11285 => x"74000000",
         11286 => x"494f4354",
         11287 => x"4c205244",
         11288 => x"20696e74",
         11289 => x"65727275",
         11290 => x"70740000",
         11291 => x"494f4354",
         11292 => x"4c205752",
         11293 => x"20696e74",
         11294 => x"65727275",
         11295 => x"70740000",
         11296 => x"55415254",
         11297 => x"30205258",
         11298 => x"20696e74",
         11299 => x"65727275",
         11300 => x"70740000",
         11301 => x"55415254",
         11302 => x"30205458",
         11303 => x"20696e74",
         11304 => x"65727275",
         11305 => x"70740000",
         11306 => x"55415254",
         11307 => x"31205258",
         11308 => x"20696e74",
         11309 => x"65727275",
         11310 => x"70740000",
         11311 => x"55415254",
         11312 => x"31205458",
         11313 => x"20696e74",
         11314 => x"65727275",
         11315 => x"70740000",
         11316 => x"53657474",
         11317 => x"696e6720",
         11318 => x"75702074",
         11319 => x"696d6572",
         11320 => x"2e2e2e00",
         11321 => x"456e6162",
         11322 => x"6c696e67",
         11323 => x"2074696d",
         11324 => x"65722e2e",
         11325 => x"2e000000",
         11326 => x"6175746f",
         11327 => x"65786563",
         11328 => x"2e626174",
         11329 => x"00000000",
         11330 => x"7a4f532e",
         11331 => x"68737400",
         11332 => x"303a0000",
         11333 => x"4661696c",
         11334 => x"65642074",
         11335 => x"6f20696e",
         11336 => x"69746961",
         11337 => x"6c697365",
         11338 => x"20736420",
         11339 => x"63617264",
         11340 => x"20302c20",
         11341 => x"706c6561",
         11342 => x"73652069",
         11343 => x"6e697420",
         11344 => x"6d616e75",
         11345 => x"616c6c79",
         11346 => x"2e000000",
         11347 => x"2a200000",
         11348 => x"436c6561",
         11349 => x"72696e67",
         11350 => x"2e2e2e2e",
         11351 => x"00000000",
         11352 => x"436f7079",
         11353 => x"696e672e",
         11354 => x"2e2e0000",
         11355 => x"436f6d70",
         11356 => x"6172696e",
         11357 => x"672e2e2e",
         11358 => x"00000000",
         11359 => x"2530386c",
         11360 => x"78282530",
         11361 => x"3878292d",
         11362 => x"3e253038",
         11363 => x"6c782825",
         11364 => x"30387829",
         11365 => x"0a000000",
         11366 => x"44756d70",
         11367 => x"204d656d",
         11368 => x"6f727900",
         11369 => x"0a436f6d",
         11370 => x"706c6574",
         11371 => x"652e0000",
         11372 => x"2530386c",
         11373 => x"58202530",
         11374 => x"32582d00",
         11375 => x"3f3f3f00",
         11376 => x"2530386c",
         11377 => x"58202530",
         11378 => x"34582d00",
         11379 => x"2530386c",
         11380 => x"58202530",
         11381 => x"386c582d",
         11382 => x"00000000",
         11383 => x"45786563",
         11384 => x"7574696e",
         11385 => x"6720636f",
         11386 => x"64652040",
         11387 => x"20253038",
         11388 => x"6c78202e",
         11389 => x"2e2e0a00",
         11390 => x"43616c6c",
         11391 => x"696e6720",
         11392 => x"636f6465",
         11393 => x"20402025",
         11394 => x"30386c78",
         11395 => x"202e2e2e",
         11396 => x"0a000000",
         11397 => x"43616c6c",
         11398 => x"20726574",
         11399 => x"75726e65",
         11400 => x"6420636f",
         11401 => x"64652028",
         11402 => x"2564292e",
         11403 => x"0a000000",
         11404 => x"52657374",
         11405 => x"61727469",
         11406 => x"6e672061",
         11407 => x"70706c69",
         11408 => x"63617469",
         11409 => x"6f6e2e2e",
         11410 => x"2e000000",
         11411 => x"436f6c64",
         11412 => x"20726562",
         11413 => x"6f6f7469",
         11414 => x"6e672e2e",
         11415 => x"2e000000",
         11416 => x"5a505500",
         11417 => x"62696e00",
         11418 => x"25643a5c",
         11419 => x"25735c25",
         11420 => x"732e2573",
         11421 => x"00000000",
         11422 => x"25643a5c",
         11423 => x"25735c25",
         11424 => x"73000000",
         11425 => x"25643a5c",
         11426 => x"25730000",
         11427 => x"42616420",
         11428 => x"636f6d6d",
         11429 => x"616e642e",
         11430 => x"00000000",
         11431 => x"52756e6e",
         11432 => x"696e672e",
         11433 => x"2e2e0000",
         11434 => x"456e6162",
         11435 => x"6c696e67",
         11436 => x"20696e74",
         11437 => x"65727275",
         11438 => x"7074732e",
         11439 => x"2e2e0000",
         11440 => x"25642f25",
         11441 => x"642f2564",
         11442 => x"2025643a",
         11443 => x"25643a25",
         11444 => x"642e2564",
         11445 => x"25640a00",
         11446 => x"536f4320",
         11447 => x"436f6e66",
         11448 => x"69677572",
         11449 => x"6174696f",
         11450 => x"6e000000",
         11451 => x"20286672",
         11452 => x"6f6d2053",
         11453 => x"6f432063",
         11454 => x"6f6e6669",
         11455 => x"67290000",
         11456 => x"3a0a4465",
         11457 => x"76696365",
         11458 => x"7320696d",
         11459 => x"706c656d",
         11460 => x"656e7465",
         11461 => x"643a0000",
         11462 => x"20202020",
         11463 => x"57422053",
         11464 => x"4452414d",
         11465 => x"20202825",
         11466 => x"3038583a",
         11467 => x"25303858",
         11468 => x"292e0a00",
         11469 => x"20202020",
         11470 => x"53445241",
         11471 => x"4d202020",
         11472 => x"20202825",
         11473 => x"3038583a",
         11474 => x"25303858",
         11475 => x"292e0a00",
         11476 => x"20202020",
         11477 => x"494e534e",
         11478 => x"20425241",
         11479 => x"4d202825",
         11480 => x"3038583a",
         11481 => x"25303858",
         11482 => x"292e0a00",
         11483 => x"20202020",
         11484 => x"4252414d",
         11485 => x"20202020",
         11486 => x"20202825",
         11487 => x"3038583a",
         11488 => x"25303858",
         11489 => x"292e0a00",
         11490 => x"20202020",
         11491 => x"52414d20",
         11492 => x"20202020",
         11493 => x"20202825",
         11494 => x"3038583a",
         11495 => x"25303858",
         11496 => x"292e0a00",
         11497 => x"20202020",
         11498 => x"53442043",
         11499 => x"41524420",
         11500 => x"20202844",
         11501 => x"65766963",
         11502 => x"6573203d",
         11503 => x"25303264",
         11504 => x"292e0a00",
         11505 => x"20202020",
         11506 => x"54494d45",
         11507 => x"52312020",
         11508 => x"20202854",
         11509 => x"696d6572",
         11510 => x"7320203d",
         11511 => x"25303264",
         11512 => x"292e0a00",
         11513 => x"20202020",
         11514 => x"494e5452",
         11515 => x"20435452",
         11516 => x"4c202843",
         11517 => x"68616e6e",
         11518 => x"656c733d",
         11519 => x"25303264",
         11520 => x"292e0a00",
         11521 => x"20202020",
         11522 => x"57495348",
         11523 => x"424f4e45",
         11524 => x"20425553",
         11525 => x"00000000",
         11526 => x"20202020",
         11527 => x"57422049",
         11528 => x"32430000",
         11529 => x"20202020",
         11530 => x"494f4354",
         11531 => x"4c000000",
         11532 => x"20202020",
         11533 => x"50533200",
         11534 => x"20202020",
         11535 => x"53504900",
         11536 => x"41646472",
         11537 => x"65737365",
         11538 => x"733a0000",
         11539 => x"20202020",
         11540 => x"43505520",
         11541 => x"52657365",
         11542 => x"74205665",
         11543 => x"63746f72",
         11544 => x"20416464",
         11545 => x"72657373",
         11546 => x"203d2025",
         11547 => x"3038580a",
         11548 => x"00000000",
         11549 => x"20202020",
         11550 => x"43505520",
         11551 => x"4d656d6f",
         11552 => x"72792053",
         11553 => x"74617274",
         11554 => x"20416464",
         11555 => x"72657373",
         11556 => x"203d2025",
         11557 => x"3038580a",
         11558 => x"00000000",
         11559 => x"20202020",
         11560 => x"53746163",
         11561 => x"6b205374",
         11562 => x"61727420",
         11563 => x"41646472",
         11564 => x"65737320",
         11565 => x"20202020",
         11566 => x"203d2025",
         11567 => x"3038580a",
         11568 => x"00000000",
         11569 => x"4d697363",
         11570 => x"3a000000",
         11571 => x"20202020",
         11572 => x"5a505520",
         11573 => x"49642020",
         11574 => x"20202020",
         11575 => x"20202020",
         11576 => x"20202020",
         11577 => x"20202020",
         11578 => x"203d2025",
         11579 => x"3034580a",
         11580 => x"00000000",
         11581 => x"20202020",
         11582 => x"53797374",
         11583 => x"656d2043",
         11584 => x"6c6f636b",
         11585 => x"20467265",
         11586 => x"71202020",
         11587 => x"20202020",
         11588 => x"203d2025",
         11589 => x"642e2530",
         11590 => x"34644d48",
         11591 => x"7a0a0000",
         11592 => x"20202020",
         11593 => x"53445241",
         11594 => x"4d20436c",
         11595 => x"6f636b20",
         11596 => x"46726571",
         11597 => x"20202020",
         11598 => x"20202020",
         11599 => x"203d2025",
         11600 => x"642e2530",
         11601 => x"34644d48",
         11602 => x"7a0a0000",
         11603 => x"20202020",
         11604 => x"57697368",
         11605 => x"626f6e65",
         11606 => x"20534452",
         11607 => x"414d2043",
         11608 => x"6c6f636b",
         11609 => x"20467265",
         11610 => x"713d2025",
         11611 => x"642e2530",
         11612 => x"34644d48",
         11613 => x"7a0a0000",
         11614 => x"536d616c",
         11615 => x"6c000000",
         11616 => x"4d656469",
         11617 => x"756d0000",
         11618 => x"466c6578",
         11619 => x"00000000",
         11620 => x"45564f00",
         11621 => x"45564f6d",
         11622 => x"00000000",
         11623 => x"556e6b6e",
         11624 => x"6f776e00",
         11625 => x"00009700",
         11626 => x"01000000",
         11627 => x"00000002",
         11628 => x"000096fc",
         11629 => x"01000000",
         11630 => x"00000003",
         11631 => x"000096f8",
         11632 => x"01000000",
         11633 => x"00000004",
         11634 => x"000096f4",
         11635 => x"01000000",
         11636 => x"00000005",
         11637 => x"000096f0",
         11638 => x"01000000",
         11639 => x"00000006",
         11640 => x"000096ec",
         11641 => x"01000000",
         11642 => x"00000007",
         11643 => x"000096e8",
         11644 => x"01000000",
         11645 => x"00000001",
         11646 => x"000096e4",
         11647 => x"01000000",
         11648 => x"00000008",
         11649 => x"000096e0",
         11650 => x"01000000",
         11651 => x"0000000b",
         11652 => x"000096dc",
         11653 => x"01000000",
         11654 => x"00000009",
         11655 => x"000096d8",
         11656 => x"01000000",
         11657 => x"0000000a",
         11658 => x"000096d4",
         11659 => x"04000000",
         11660 => x"0000000d",
         11661 => x"000096d0",
         11662 => x"04000000",
         11663 => x"0000000c",
         11664 => x"000096cc",
         11665 => x"04000000",
         11666 => x"0000000e",
         11667 => x"000096c8",
         11668 => x"03000000",
         11669 => x"0000000f",
         11670 => x"000096c4",
         11671 => x"04000000",
         11672 => x"0000000f",
         11673 => x"000096c0",
         11674 => x"04000000",
         11675 => x"00000010",
         11676 => x"000096bc",
         11677 => x"04000000",
         11678 => x"00000011",
         11679 => x"000096b8",
         11680 => x"03000000",
         11681 => x"00000012",
         11682 => x"000096b4",
         11683 => x"03000000",
         11684 => x"00000013",
         11685 => x"000096b0",
         11686 => x"03000000",
         11687 => x"00000014",
         11688 => x"000096ac",
         11689 => x"03000000",
         11690 => x"00000015",
         11691 => x"1b5b4400",
         11692 => x"1b5b4300",
         11693 => x"1b5b4200",
         11694 => x"1b5b4100",
         11695 => x"1b5b367e",
         11696 => x"1b5b357e",
         11697 => x"1b5b347e",
         11698 => x"1b304600",
         11699 => x"1b5b337e",
         11700 => x"1b5b327e",
         11701 => x"1b5b317e",
         11702 => x"10000000",
         11703 => x"0e000000",
         11704 => x"0d000000",
         11705 => x"0b000000",
         11706 => x"08000000",
         11707 => x"06000000",
         11708 => x"05000000",
         11709 => x"04000000",
         11710 => x"03000000",
         11711 => x"02000000",
         11712 => x"01000000",
         11713 => x"68697374",
         11714 => x"6f727900",
         11715 => x"68697374",
         11716 => x"00000000",
         11717 => x"21000000",
         11718 => x"2530346c",
         11719 => x"75202025",
         11720 => x"730a0000",
         11721 => x"4661696c",
         11722 => x"65642074",
         11723 => x"6f207265",
         11724 => x"73657420",
         11725 => x"74686520",
         11726 => x"68697374",
         11727 => x"6f727920",
         11728 => x"66696c65",
         11729 => x"20746f20",
         11730 => x"454f462e",
         11731 => x"00000000",
         11732 => x"43616e6e",
         11733 => x"6f74206f",
         11734 => x"70656e2f",
         11735 => x"63726561",
         11736 => x"74652068",
         11737 => x"6973746f",
         11738 => x"72792066",
         11739 => x"696c652c",
         11740 => x"20646973",
         11741 => x"61626c69",
         11742 => x"6e672e00",
         11743 => x"53440000",
         11744 => x"222a2b2c",
         11745 => x"3a3b3c3d",
         11746 => x"3e3f5b5d",
         11747 => x"7c7f0000",
         11748 => x"46415400",
         11749 => x"46415433",
         11750 => x"32000000",
         11751 => x"ebfe904d",
         11752 => x"53444f53",
         11753 => x"352e3000",
         11754 => x"4e4f204e",
         11755 => x"414d4520",
         11756 => x"20202046",
         11757 => x"41543332",
         11758 => x"20202000",
         11759 => x"4e4f204e",
         11760 => x"414d4520",
         11761 => x"20202046",
         11762 => x"41542020",
         11763 => x"20202000",
         11764 => x"0000977c",
         11765 => x"00000000",
         11766 => x"00000000",
         11767 => x"00000000",
         11768 => x"809a4541",
         11769 => x"8e418f80",
         11770 => x"45454549",
         11771 => x"49498e8f",
         11772 => x"9092924f",
         11773 => x"994f5555",
         11774 => x"59999a9b",
         11775 => x"9c9d9e9f",
         11776 => x"41494f55",
         11777 => x"a5a5a6a7",
         11778 => x"a8a9aaab",
         11779 => x"acadaeaf",
         11780 => x"b0b1b2b3",
         11781 => x"b4b5b6b7",
         11782 => x"b8b9babb",
         11783 => x"bcbdbebf",
         11784 => x"c0c1c2c3",
         11785 => x"c4c5c6c7",
         11786 => x"c8c9cacb",
         11787 => x"cccdcecf",
         11788 => x"d0d1d2d3",
         11789 => x"d4d5d6d7",
         11790 => x"d8d9dadb",
         11791 => x"dcdddedf",
         11792 => x"e0e1e2e3",
         11793 => x"e4e5e6e7",
         11794 => x"e8e9eaeb",
         11795 => x"ecedeeef",
         11796 => x"f0f1f2f3",
         11797 => x"f4f5f6f7",
         11798 => x"f8f9fafb",
         11799 => x"fcfdfeff",
         11800 => x"2b2e2c3b",
         11801 => x"3d5b5d2f",
         11802 => x"5c222a3a",
         11803 => x"3c3e3f7c",
         11804 => x"7f000000",
         11805 => x"00010004",
         11806 => x"00100040",
         11807 => x"01000200",
         11808 => x"00000000",
         11809 => x"00010002",
         11810 => x"00040008",
         11811 => x"00100020",
         11812 => x"00000000",
         11813 => x"00000000",
         11814 => x"00008cec",
         11815 => x"01020100",
         11816 => x"00000000",
         11817 => x"00000000",
         11818 => x"00008cf4",
         11819 => x"01040100",
         11820 => x"00000000",
         11821 => x"00000000",
         11822 => x"00008cfc",
         11823 => x"01140300",
         11824 => x"00000000",
         11825 => x"00000000",
         11826 => x"00008d04",
         11827 => x"012b0300",
         11828 => x"00000000",
         11829 => x"00000000",
         11830 => x"00008d0c",
         11831 => x"01300300",
         11832 => x"00000000",
         11833 => x"00000000",
         11834 => x"00008d14",
         11835 => x"013c0400",
         11836 => x"00000000",
         11837 => x"00000000",
         11838 => x"00008d1c",
         11839 => x"013d0400",
         11840 => x"00000000",
         11841 => x"00000000",
         11842 => x"00008d24",
         11843 => x"013f0400",
         11844 => x"00000000",
         11845 => x"00000000",
         11846 => x"00008d2c",
         11847 => x"01400400",
         11848 => x"00000000",
         11849 => x"00000000",
         11850 => x"00008d34",
         11851 => x"01410400",
         11852 => x"00000000",
         11853 => x"00000000",
         11854 => x"00008d38",
         11855 => x"01420400",
         11856 => x"00000000",
         11857 => x"00000000",
         11858 => x"00008d3c",
         11859 => x"01430400",
         11860 => x"00000000",
         11861 => x"00000000",
         11862 => x"00008d40",
         11863 => x"01500500",
         11864 => x"00000000",
         11865 => x"00000000",
         11866 => x"00008d44",
         11867 => x"01510500",
         11868 => x"00000000",
         11869 => x"00000000",
         11870 => x"00008d48",
         11871 => x"01540500",
         11872 => x"00000000",
         11873 => x"00000000",
         11874 => x"00008d4c",
         11875 => x"01550500",
         11876 => x"00000000",
         11877 => x"00000000",
         11878 => x"00008d50",
         11879 => x"01790700",
         11880 => x"00000000",
         11881 => x"00000000",
         11882 => x"00008d58",
         11883 => x"01780700",
         11884 => x"00000000",
         11885 => x"00000000",
         11886 => x"00008d5c",
         11887 => x"01820800",
         11888 => x"00000000",
         11889 => x"00000000",
         11890 => x"00008d64",
         11891 => x"01830800",
         11892 => x"00000000",
         11893 => x"00000000",
         11894 => x"00008d6c",
         11895 => x"01850800",
         11896 => x"00000000",
         11897 => x"00000000",
         11898 => x"00008d74",
         11899 => x"01870800",
         11900 => x"00000000",
         11901 => x"00000000",
         11902 => x"00008d7c",
         11903 => x"018c0900",
         11904 => x"00000000",
         11905 => x"00000000",
         11906 => x"00008d84",
         11907 => x"018d0900",
         11908 => x"00000000",
         11909 => x"00000000",
         11910 => x"00008d8c",
         11911 => x"018e0900",
         11912 => x"00000000",
         11913 => x"00000000",
         11914 => x"00008d94",
         11915 => x"018f0900",
         11916 => x"00000000",
         11917 => x"00000000",
         11918 => x"00000000",
         11919 => x"00000000",
         11920 => x"00007fff",
         11921 => x"00000000",
         11922 => x"00007fff",
         11923 => x"00010000",
         11924 => x"00007fff",
         11925 => x"00010000",
         11926 => x"00810000",
         11927 => x"01000000",
         11928 => x"017fffff",
         11929 => x"00000000",
         11930 => x"00000000",
         11931 => x"00007800",
         11932 => x"00000000",
         11933 => x"05f5e100",
         11934 => x"05f5e100",
         11935 => x"05f5e100",
         11936 => x"00000000",
         11937 => x"01010101",
         11938 => x"01010101",
         11939 => x"01011001",
         11940 => x"01000000",
         11941 => x"00000000",
         11942 => x"00000000",
         11943 => x"00000000",
         11944 => x"00000000",
         11945 => x"00000000",
         11946 => x"00000000",
         11947 => x"00000000",
         11948 => x"00000000",
         11949 => x"00000000",
         11950 => x"00000000",
         11951 => x"00000000",
         11952 => x"00000000",
         11953 => x"00000000",
         11954 => x"00000000",
         11955 => x"00000000",
         11956 => x"00000000",
         11957 => x"00000000",
         11958 => x"00000000",
         11959 => x"00000000",
         11960 => x"00000000",
         11961 => x"00000000",
         11962 => x"00000000",
         11963 => x"00000000",
         11964 => x"00000000",
         11965 => x"00009704",
         11966 => x"01000000",
         11967 => x"0000970c",
         11968 => x"01000000",
         11969 => x"00009714",
         11970 => x"02000000",
         11971 => x"00000000",
         11972 => x"00000000",
         11973 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

