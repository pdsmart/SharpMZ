-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b83ff",
             1 => x"f80d0b0b",
             2 => x"0b939b04",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b92",
            73 => x"ff040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b92e2",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b81e7",
           162 => x"fc738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"92e70400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b99",
           171 => x"fb2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b9b",
           179 => x"e72d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"95040b0b",
           269 => x"0b8ca504",
           270 => x"0b0b0b8c",
           271 => x"b5040b0b",
           272 => x"0b8cc504",
           273 => x"0b0b0b8c",
           274 => x"d5040b0b",
           275 => x"0b8ce504",
           276 => x"0b0b0b8c",
           277 => x"f5040b0b",
           278 => x"0b8d8504",
           279 => x"0b0b0b8d",
           280 => x"95040b0b",
           281 => x"0b8da504",
           282 => x"0b0b0b8d",
           283 => x"b5040b0b",
           284 => x"0b8dc504",
           285 => x"0b0b0b8d",
           286 => x"d5040b0b",
           287 => x"0b8de504",
           288 => x"0b0b0b8d",
           289 => x"f5040b0b",
           290 => x"0b8e8404",
           291 => x"0b0b0b8e",
           292 => x"93040b0b",
           293 => x"0b8ea204",
           294 => x"0b0b0b8e",
           295 => x"b2040b0b",
           296 => x"0b8ec204",
           297 => x"0b0b0b8e",
           298 => x"d2040b0b",
           299 => x"0b8ee204",
           300 => x"0b0b0b8e",
           301 => x"f2040b0b",
           302 => x"0b8f8204",
           303 => x"0b0b0b8f",
           304 => x"92040b0b",
           305 => x"0b8fa204",
           306 => x"0b0b0b8f",
           307 => x"b2040b0b",
           308 => x"0b8fc204",
           309 => x"0b0b0b8f",
           310 => x"d2040b0b",
           311 => x"0b8fe204",
           312 => x"0b0b0b8f",
           313 => x"f2040b0b",
           314 => x"0b908204",
           315 => x"0b0b0b90",
           316 => x"92040b0b",
           317 => x"0b90a204",
           318 => x"0b0b0b90",
           319 => x"b2040b0b",
           320 => x"0b90c204",
           321 => x"0b0b0b90",
           322 => x"d2040b0b",
           323 => x"0b90e204",
           324 => x"0b0b0b90",
           325 => x"f2040b0b",
           326 => x"0b918204",
           327 => x"0b0b0b91",
           328 => x"92040b0b",
           329 => x"0b91a204",
           330 => x"0b0b0b91",
           331 => x"b2040b0b",
           332 => x"0b91c204",
           333 => x"0b0b0b91",
           334 => x"d2040b0b",
           335 => x"0b91e204",
           336 => x"0b0b0b91",
           337 => x"f2040b0b",
           338 => x"0b928204",
           339 => x"0b0b0b92",
           340 => x"91040b0b",
           341 => x"0b92a004",
           342 => x"0b0b0b92",
           343 => x"b004ffff",
           344 => x"ffffffff",
           345 => x"ffffffff",
           346 => x"ffffffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"048285f8",
           386 => x"0c80c18c",
           387 => x"2d8285f8",
           388 => x"0882a090",
           389 => x"048285f8",
           390 => x"0c80ce8e",
           391 => x"2d8285f8",
           392 => x"0882a090",
           393 => x"048285f8",
           394 => x"0c80cecd",
           395 => x"2d8285f8",
           396 => x"0882a090",
           397 => x"048285f8",
           398 => x"0c80ceeb",
           399 => x"2d8285f8",
           400 => x"0882a090",
           401 => x"048285f8",
           402 => x"0c80d5b5",
           403 => x"2d8285f8",
           404 => x"0882a090",
           405 => x"048285f8",
           406 => x"0c80d6b6",
           407 => x"2d8285f8",
           408 => x"0882a090",
           409 => x"048285f8",
           410 => x"0c80cf8e",
           411 => x"2d8285f8",
           412 => x"0882a090",
           413 => x"048285f8",
           414 => x"0c80d6d3",
           415 => x"2d8285f8",
           416 => x"0882a090",
           417 => x"048285f8",
           418 => x"0c80d8cf",
           419 => x"2d8285f8",
           420 => x"0882a090",
           421 => x"048285f8",
           422 => x"0c80d4db",
           423 => x"2d8285f8",
           424 => x"0882a090",
           425 => x"048285f8",
           426 => x"0c80cfc0",
           427 => x"2d8285f8",
           428 => x"0882a090",
           429 => x"048285f8",
           430 => x"0c80d4f1",
           431 => x"2d8285f8",
           432 => x"0882a090",
           433 => x"048285f8",
           434 => x"0c80d595",
           435 => x"2d8285f8",
           436 => x"0882a090",
           437 => x"048285f8",
           438 => x"0c80c395",
           439 => x"2d8285f8",
           440 => x"0882a090",
           441 => x"048285f8",
           442 => x"0c80c3e4",
           443 => x"2d8285f8",
           444 => x"0882a090",
           445 => x"048285f8",
           446 => x"0cbbc42d",
           447 => x"8285f808",
           448 => x"82a09004",
           449 => x"8285f80c",
           450 => x"bdbd2d82",
           451 => x"85f80882",
           452 => x"a0900482",
           453 => x"85f80cbe",
           454 => x"f02d8285",
           455 => x"f80882a0",
           456 => x"90048285",
           457 => x"f80c81aa",
           458 => x"bc2d8285",
           459 => x"f80882a0",
           460 => x"90048285",
           461 => x"f80c81b7",
           462 => x"af2d8285",
           463 => x"f80882a0",
           464 => x"90048285",
           465 => x"f80c81af",
           466 => x"a32d8285",
           467 => x"f80882a0",
           468 => x"90048285",
           469 => x"f80c81b2",
           470 => x"a02d8285",
           471 => x"f80882a0",
           472 => x"90048285",
           473 => x"f80c81bc",
           474 => x"bd2d8285",
           475 => x"f80882a0",
           476 => x"90048285",
           477 => x"f80c81c5",
           478 => x"a82d8285",
           479 => x"f80882a0",
           480 => x"90048285",
           481 => x"f80c81b6",
           482 => x"912d8285",
           483 => x"f80882a0",
           484 => x"90048285",
           485 => x"f80c81bf",
           486 => x"de2d8285",
           487 => x"f80882a0",
           488 => x"90048285",
           489 => x"f80c81c0",
           490 => x"fd2d8285",
           491 => x"f80882a0",
           492 => x"90048285",
           493 => x"f80c81c1",
           494 => x"9c2d8285",
           495 => x"f80882a0",
           496 => x"90048285",
           497 => x"f80c81c9",
           498 => x"912d8285",
           499 => x"f80882a0",
           500 => x"90048285",
           501 => x"f80c81c6",
           502 => x"f52d8285",
           503 => x"f80882a0",
           504 => x"90048285",
           505 => x"f80c81cb",
           506 => x"e52d8285",
           507 => x"f80882a0",
           508 => x"90048285",
           509 => x"f80c81c2",
           510 => x"a22d8285",
           511 => x"f80882a0",
           512 => x"90048285",
           513 => x"f80c81ce",
           514 => x"e52d8285",
           515 => x"f80882a0",
           516 => x"90048285",
           517 => x"f80c81cf",
           518 => x"e62d8285",
           519 => x"f80882a0",
           520 => x"90048285",
           521 => x"f80c81b8",
           522 => x"8f2d8285",
           523 => x"f80882a0",
           524 => x"90048285",
           525 => x"f80c81b7",
           526 => x"e82d8285",
           527 => x"f80882a0",
           528 => x"90048285",
           529 => x"f80c81b9",
           530 => x"932d8285",
           531 => x"f80882a0",
           532 => x"90048285",
           533 => x"f80c81c2",
           534 => x"f92d8285",
           535 => x"f80882a0",
           536 => x"90048285",
           537 => x"f80c81d0",
           538 => x"d72d8285",
           539 => x"f80882a0",
           540 => x"90048285",
           541 => x"f80c81d2",
           542 => x"e52d8285",
           543 => x"f80882a0",
           544 => x"90048285",
           545 => x"f80c81d6",
           546 => x"a72d8285",
           547 => x"f80882a0",
           548 => x"90048285",
           549 => x"f80c81a9",
           550 => x"db2d8285",
           551 => x"f80882a0",
           552 => x"90048285",
           553 => x"f80c81d9",
           554 => x"952d8285",
           555 => x"f80882a0",
           556 => x"90048285",
           557 => x"f80c81e7",
           558 => x"d92d8285",
           559 => x"f80882a0",
           560 => x"90048285",
           561 => x"f80c81e5",
           562 => x"c02d8285",
           563 => x"f80882a0",
           564 => x"90048285",
           565 => x"f80c80fa",
           566 => x"e82d8285",
           567 => x"f80882a0",
           568 => x"90048285",
           569 => x"f80c80fc",
           570 => x"d22d8285",
           571 => x"f80882a0",
           572 => x"90048285",
           573 => x"f80c80fe",
           574 => x"b62d8285",
           575 => x"f80882a0",
           576 => x"90048285",
           577 => x"f80cbbed",
           578 => x"2d8285f8",
           579 => x"0882a090",
           580 => x"048285f8",
           581 => x"0cbd932d",
           582 => x"8285f808",
           583 => x"82a09004",
           584 => x"8285f80c",
           585 => x"80c0802d",
           586 => x"8285f808",
           587 => x"82a09004",
           588 => x"8285f80c",
           589 => x"a1fd2d82",
           590 => x"85f80882",
           591 => x"a090043c",
           592 => x"04000010",
           593 => x"10101010",
           594 => x"10101010",
           595 => x"10101010",
           596 => x"10101010",
           597 => x"10101010",
           598 => x"10101010",
           599 => x"10101010",
           600 => x"10105351",
           601 => x"04000073",
           602 => x"81ff0673",
           603 => x"83060981",
           604 => x"05830510",
           605 => x"10102b07",
           606 => x"72fc060c",
           607 => x"51510472",
           608 => x"72807281",
           609 => x"06ff0509",
           610 => x"72060571",
           611 => x"1052720a",
           612 => x"100a5372",
           613 => x"ed385151",
           614 => x"53510482",
           615 => x"85ec7082",
           616 => x"9da8278e",
           617 => x"38807170",
           618 => x"8405530c",
           619 => x"0b0b0b93",
           620 => x"9e048c81",
           621 => x"51ba9d04",
           622 => x"008285f8",
           623 => x"08028285",
           624 => x"f80cfe3d",
           625 => x"0d8285f8",
           626 => x"08880508",
           627 => x"8285f808",
           628 => x"fc050c82",
           629 => x"85f808fc",
           630 => x"05085271",
           631 => x"338285f8",
           632 => x"08fc0508",
           633 => x"81058285",
           634 => x"f808fc05",
           635 => x"0c7081ff",
           636 => x"06515170",
           637 => x"802e8338",
           638 => x"da398285",
           639 => x"f808fc05",
           640 => x"08ff0582",
           641 => x"85f808fc",
           642 => x"050c8285",
           643 => x"f808fc05",
           644 => x"088285f8",
           645 => x"08880508",
           646 => x"31708285",
           647 => x"ec0c5184",
           648 => x"3d0d8285",
           649 => x"f80c0482",
           650 => x"85f80802",
           651 => x"8285f80c",
           652 => x"fe3d0d82",
           653 => x"85f80888",
           654 => x"05088285",
           655 => x"f808fc05",
           656 => x"0c8285f8",
           657 => x"088c0508",
           658 => x"52713382",
           659 => x"85f8088c",
           660 => x"05088105",
           661 => x"8285f808",
           662 => x"8c050c82",
           663 => x"85f808fc",
           664 => x"05085351",
           665 => x"70723482",
           666 => x"85f808fc",
           667 => x"05088105",
           668 => x"8285f808",
           669 => x"fc050c70",
           670 => x"81ff0651",
           671 => x"70802e84",
           672 => x"38ffbe39",
           673 => x"8285f808",
           674 => x"88050870",
           675 => x"8285ec0c",
           676 => x"51843d0d",
           677 => x"8285f80c",
           678 => x"048285f8",
           679 => x"08028285",
           680 => x"f80cfd3d",
           681 => x"0d8285f8",
           682 => x"08880508",
           683 => x"8285f808",
           684 => x"fc050c82",
           685 => x"85f8088c",
           686 => x"05088285",
           687 => x"f808f805",
           688 => x"0c8285f8",
           689 => x"08900508",
           690 => x"802e80e5",
           691 => x"388285f8",
           692 => x"08900508",
           693 => x"81058285",
           694 => x"f8089005",
           695 => x"0c8285f8",
           696 => x"08900508",
           697 => x"ff058285",
           698 => x"f8089005",
           699 => x"0c8285f8",
           700 => x"08900508",
           701 => x"802eba38",
           702 => x"8285f808",
           703 => x"f8050851",
           704 => x"70338285",
           705 => x"f808f805",
           706 => x"08810582",
           707 => x"85f808f8",
           708 => x"050c8285",
           709 => x"f808fc05",
           710 => x"08525271",
           711 => x"71348285",
           712 => x"f808fc05",
           713 => x"08810582",
           714 => x"85f808fc",
           715 => x"050cffad",
           716 => x"398285f8",
           717 => x"08880508",
           718 => x"708285ec",
           719 => x"0c51853d",
           720 => x"0d8285f8",
           721 => x"0c048285",
           722 => x"f8080282",
           723 => x"85f80cfd",
           724 => x"3d0d8285",
           725 => x"f8089005",
           726 => x"08802e81",
           727 => x"f4388285",
           728 => x"f8088c05",
           729 => x"08527133",
           730 => x"8285f808",
           731 => x"8c050881",
           732 => x"058285f8",
           733 => x"088c050c",
           734 => x"8285f808",
           735 => x"88050870",
           736 => x"337281ff",
           737 => x"06535454",
           738 => x"5171712e",
           739 => x"843880ce",
           740 => x"398285f8",
           741 => x"08880508",
           742 => x"52713382",
           743 => x"85f80888",
           744 => x"05088105",
           745 => x"8285f808",
           746 => x"88050c70",
           747 => x"81ff0651",
           748 => x"51708d38",
           749 => x"800b8285",
           750 => x"f808fc05",
           751 => x"0c819b39",
           752 => x"8285f808",
           753 => x"900508ff",
           754 => x"058285f8",
           755 => x"0890050c",
           756 => x"8285f808",
           757 => x"90050880",
           758 => x"2e8438ff",
           759 => x"81398285",
           760 => x"f8089005",
           761 => x"08802e80",
           762 => x"e8388285",
           763 => x"f8088805",
           764 => x"08703352",
           765 => x"53708d38",
           766 => x"ff0b8285",
           767 => x"f808fc05",
           768 => x"0c80d739",
           769 => x"8285f808",
           770 => x"8c0508ff",
           771 => x"058285f8",
           772 => x"088c050c",
           773 => x"8285f808",
           774 => x"8c050870",
           775 => x"33525270",
           776 => x"8c38810b",
           777 => x"8285f808",
           778 => x"fc050cae",
           779 => x"398285f8",
           780 => x"08880508",
           781 => x"70338285",
           782 => x"f8088c05",
           783 => x"08703372",
           784 => x"71317082",
           785 => x"85f808fc",
           786 => x"050c5355",
           787 => x"5252538a",
           788 => x"39800b82",
           789 => x"85f808fc",
           790 => x"050c8285",
           791 => x"f808fc05",
           792 => x"088285ec",
           793 => x"0c853d0d",
           794 => x"8285f80c",
           795 => x"048285f8",
           796 => x"08028285",
           797 => x"f80cfe3d",
           798 => x"0d8285f8",
           799 => x"08880508",
           800 => x"8285f808",
           801 => x"fc050c82",
           802 => x"85f80890",
           803 => x"0508802e",
           804 => x"80d43882",
           805 => x"85f80890",
           806 => x"05088105",
           807 => x"8285f808",
           808 => x"90050c82",
           809 => x"85f80890",
           810 => x"0508ff05",
           811 => x"8285f808",
           812 => x"90050c82",
           813 => x"85f80890",
           814 => x"0508802e",
           815 => x"a9388285",
           816 => x"f8088c05",
           817 => x"08517082",
           818 => x"85f808fc",
           819 => x"05085252",
           820 => x"71713482",
           821 => x"85f808fc",
           822 => x"05088105",
           823 => x"8285f808",
           824 => x"fc050cff",
           825 => x"be398285",
           826 => x"f8088805",
           827 => x"08708285",
           828 => x"ec0c5184",
           829 => x"3d0d8285",
           830 => x"f80c0482",
           831 => x"85f80802",
           832 => x"8285f80c",
           833 => x"f93d0d80",
           834 => x"0b8285f8",
           835 => x"08fc050c",
           836 => x"8285f808",
           837 => x"88050880",
           838 => x"25b93882",
           839 => x"85f80888",
           840 => x"05083082",
           841 => x"85f80888",
           842 => x"050c800b",
           843 => x"8285f808",
           844 => x"f4050c82",
           845 => x"85f808fc",
           846 => x"05088a38",
           847 => x"810b8285",
           848 => x"f808f405",
           849 => x"0c8285f8",
           850 => x"08f40508",
           851 => x"8285f808",
           852 => x"fc050c82",
           853 => x"85f8088c",
           854 => x"05088025",
           855 => x"b9388285",
           856 => x"f8088c05",
           857 => x"08308285",
           858 => x"f8088c05",
           859 => x"0c800b82",
           860 => x"85f808f0",
           861 => x"050c8285",
           862 => x"f808fc05",
           863 => x"088a3881",
           864 => x"0b8285f8",
           865 => x"08f0050c",
           866 => x"8285f808",
           867 => x"f0050882",
           868 => x"85f808fc",
           869 => x"050c8053",
           870 => x"8285f808",
           871 => x"8c050852",
           872 => x"8285f808",
           873 => x"88050851",
           874 => x"83c53f82",
           875 => x"85ec0870",
           876 => x"8285f808",
           877 => x"f8050c54",
           878 => x"8285f808",
           879 => x"fc050880",
           880 => x"2e903882",
           881 => x"85f808f8",
           882 => x"05083082",
           883 => x"85f808f8",
           884 => x"050c8285",
           885 => x"f808f805",
           886 => x"08708285",
           887 => x"ec0c5489",
           888 => x"3d0d8285",
           889 => x"f80c0482",
           890 => x"85f80802",
           891 => x"8285f80c",
           892 => x"fb3d0d80",
           893 => x"0b8285f8",
           894 => x"08fc050c",
           895 => x"8285f808",
           896 => x"88050880",
           897 => x"25993882",
           898 => x"85f80888",
           899 => x"05083082",
           900 => x"85f80888",
           901 => x"050c810b",
           902 => x"8285f808",
           903 => x"fc050c82",
           904 => x"85f8088c",
           905 => x"05088025",
           906 => x"90388285",
           907 => x"f8088c05",
           908 => x"08308285",
           909 => x"f8088c05",
           910 => x"0c815382",
           911 => x"85f8088c",
           912 => x"05085282",
           913 => x"85f80888",
           914 => x"05085182",
           915 => x"a23f8285",
           916 => x"ec087082",
           917 => x"85f808f8",
           918 => x"050c5482",
           919 => x"85f808fc",
           920 => x"0508802e",
           921 => x"90388285",
           922 => x"f808f805",
           923 => x"08308285",
           924 => x"f808f805",
           925 => x"0c8285f8",
           926 => x"08f80508",
           927 => x"708285ec",
           928 => x"0c54873d",
           929 => x"0d8285f8",
           930 => x"0c048285",
           931 => x"f8080282",
           932 => x"85f80cff",
           933 => x"3d0d800b",
           934 => x"8285f808",
           935 => x"fc050c82",
           936 => x"85f80888",
           937 => x"05088106",
           938 => x"ff117009",
           939 => x"708285f8",
           940 => x"088c0508",
           941 => x"068285f8",
           942 => x"08fc0508",
           943 => x"118285f8",
           944 => x"08fc050c",
           945 => x"8285f808",
           946 => x"88050881",
           947 => x"2a8285f8",
           948 => x"0888050c",
           949 => x"8285f808",
           950 => x"8c050810",
           951 => x"8285f808",
           952 => x"8c050c51",
           953 => x"51515182",
           954 => x"85f80888",
           955 => x"0508802e",
           956 => x"8438ffab",
           957 => x"398285f8",
           958 => x"08fc0508",
           959 => x"708285ec",
           960 => x"0c51833d",
           961 => x"0d8285f8",
           962 => x"0c048285",
           963 => x"f8080282",
           964 => x"85f80cfd",
           965 => x"3d0d8053",
           966 => x"8285f808",
           967 => x"8c050852",
           968 => x"8285f808",
           969 => x"88050851",
           970 => x"80c53f82",
           971 => x"85ec0870",
           972 => x"8285ec0c",
           973 => x"54853d0d",
           974 => x"8285f80c",
           975 => x"048285f8",
           976 => x"08028285",
           977 => x"f80cfd3d",
           978 => x"0d815382",
           979 => x"85f8088c",
           980 => x"05085282",
           981 => x"85f80888",
           982 => x"05085193",
           983 => x"3f8285ec",
           984 => x"08708285",
           985 => x"ec0c5485",
           986 => x"3d0d8285",
           987 => x"f80c0482",
           988 => x"85f80802",
           989 => x"8285f80c",
           990 => x"fd3d0d81",
           991 => x"0b8285f8",
           992 => x"08fc050c",
           993 => x"800b8285",
           994 => x"f808f805",
           995 => x"0c8285f8",
           996 => x"088c0508",
           997 => x"8285f808",
           998 => x"88050827",
           999 => x"b9388285",
          1000 => x"f808fc05",
          1001 => x"08802eae",
          1002 => x"38800b82",
          1003 => x"85f8088c",
          1004 => x"050824a2",
          1005 => x"388285f8",
          1006 => x"088c0508",
          1007 => x"108285f8",
          1008 => x"088c050c",
          1009 => x"8285f808",
          1010 => x"fc050810",
          1011 => x"8285f808",
          1012 => x"fc050cff",
          1013 => x"b8398285",
          1014 => x"f808fc05",
          1015 => x"08802e80",
          1016 => x"e1388285",
          1017 => x"f8088c05",
          1018 => x"088285f8",
          1019 => x"08880508",
          1020 => x"26ad3882",
          1021 => x"85f80888",
          1022 => x"05088285",
          1023 => x"f8088c05",
          1024 => x"08318285",
          1025 => x"f8088805",
          1026 => x"0c8285f8",
          1027 => x"08f80508",
          1028 => x"8285f808",
          1029 => x"fc050807",
          1030 => x"8285f808",
          1031 => x"f8050c82",
          1032 => x"85f808fc",
          1033 => x"0508812a",
          1034 => x"8285f808",
          1035 => x"fc050c82",
          1036 => x"85f8088c",
          1037 => x"0508812a",
          1038 => x"8285f808",
          1039 => x"8c050cff",
          1040 => x"95398285",
          1041 => x"f8089005",
          1042 => x"08802e93",
          1043 => x"388285f8",
          1044 => x"08880508",
          1045 => x"708285f8",
          1046 => x"08f4050c",
          1047 => x"51913982",
          1048 => x"85f808f8",
          1049 => x"05087082",
          1050 => x"85f808f4",
          1051 => x"050c5182",
          1052 => x"85f808f4",
          1053 => x"05088285",
          1054 => x"ec0c853d",
          1055 => x"0d8285f8",
          1056 => x"0c04f93d",
          1057 => x"0d797008",
          1058 => x"70565658",
          1059 => x"74802e80",
          1060 => x"e3389539",
          1061 => x"750851f2",
          1062 => x"a03f8285",
          1063 => x"ec081578",
          1064 => x"0c851633",
          1065 => x"5480cd39",
          1066 => x"74335473",
          1067 => x"a02e0981",
          1068 => x"06863881",
          1069 => x"1555f139",
          1070 => x"80577684",
          1071 => x"2b8280ec",
          1072 => x"05700852",
          1073 => x"56f1f23f",
          1074 => x"8285ec08",
          1075 => x"53745275",
          1076 => x"0851f4f2",
          1077 => x"3f8285ec",
          1078 => x"088b3884",
          1079 => x"16335473",
          1080 => x"812effb0",
          1081 => x"38811770",
          1082 => x"81ff0658",
          1083 => x"54997727",
          1084 => x"c938ff54",
          1085 => x"738285ec",
          1086 => x"0c893d0d",
          1087 => x"04ff3d0d",
          1088 => x"73527193",
          1089 => x"26818d38",
          1090 => x"71822b52",
          1091 => x"81e88c12",
          1092 => x"080481ea",
          1093 => x"f4518180",
          1094 => x"3981eb80",
          1095 => x"5180f939",
          1096 => x"81eb9451",
          1097 => x"80f23981",
          1098 => x"eba85180",
          1099 => x"eb3981eb",
          1100 => x"b85180e4",
          1101 => x"3981ebc8",
          1102 => x"5180dd39",
          1103 => x"81ebdc51",
          1104 => x"80d63981",
          1105 => x"ebec5180",
          1106 => x"cf3981ec",
          1107 => x"845180c8",
          1108 => x"3981ec9c",
          1109 => x"5180c139",
          1110 => x"81ecb451",
          1111 => x"bb3981ec",
          1112 => x"d051b539",
          1113 => x"81ece451",
          1114 => x"af3981ed",
          1115 => x"9051a939",
          1116 => x"81eda451",
          1117 => x"a33981ed",
          1118 => x"c4519d39",
          1119 => x"81edd851",
          1120 => x"973981ed",
          1121 => x"f0519139",
          1122 => x"81ee8851",
          1123 => x"8b3981ee",
          1124 => x"a0518539",
          1125 => x"81eeac51",
          1126 => x"abd13f83",
          1127 => x"3d0d04fb",
          1128 => x"3d0d7779",
          1129 => x"56567487",
          1130 => x"e7269238",
          1131 => x"87e85275",
          1132 => x"51f9d73f",
          1133 => x"74528285",
          1134 => x"ec085190",
          1135 => x"3987e852",
          1136 => x"7451fac6",
          1137 => x"3f8285ec",
          1138 => x"08527551",
          1139 => x"fabc3f82",
          1140 => x"85ec0854",
          1141 => x"79537552",
          1142 => x"81eebc51",
          1143 => x"b0fd3f87",
          1144 => x"3d0d04ec",
          1145 => x"3d0d6602",
          1146 => x"840580e3",
          1147 => x"05335b57",
          1148 => x"80687809",
          1149 => x"8105707a",
          1150 => x"07732551",
          1151 => x"57595978",
          1152 => x"567787ff",
          1153 => x"26833881",
          1154 => x"56747607",
          1155 => x"7081ff06",
          1156 => x"51559356",
          1157 => x"74818638",
          1158 => x"81537652",
          1159 => x"8c3d7052",
          1160 => x"56818698",
          1161 => x"3f8285ec",
          1162 => x"08578285",
          1163 => x"ec08b938",
          1164 => x"8285ec08",
          1165 => x"87c09888",
          1166 => x"0c8285ec",
          1167 => x"0859963d",
          1168 => x"d4055484",
          1169 => x"80537752",
          1170 => x"7551818a",
          1171 => x"d63f8285",
          1172 => x"ec085782",
          1173 => x"85ec0890",
          1174 => x"387a5574",
          1175 => x"802e8938",
          1176 => x"74197519",
          1177 => x"5959d739",
          1178 => x"963dd805",
          1179 => x"518192bf",
          1180 => x"3f760981",
          1181 => x"05707807",
          1182 => x"80257b09",
          1183 => x"8105709f",
          1184 => x"2a720651",
          1185 => x"57515674",
          1186 => x"802e9038",
          1187 => x"81eee053",
          1188 => x"87c09888",
          1189 => x"08527851",
          1190 => x"fe853f76",
          1191 => x"56758285",
          1192 => x"ec0c963d",
          1193 => x"0d04f93d",
          1194 => x"0d7b0284",
          1195 => x"05b30533",
          1196 => x"5758ff57",
          1197 => x"80537a52",
          1198 => x"7951fea7",
          1199 => x"3f8285ec",
          1200 => x"08a43875",
          1201 => x"802e8838",
          1202 => x"75812e98",
          1203 => x"38983960",
          1204 => x"557f5482",
          1205 => x"85ec537e",
          1206 => x"527d5177",
          1207 => x"2d8285ec",
          1208 => x"08578339",
          1209 => x"77047682",
          1210 => x"85ec0c89",
          1211 => x"3d0d04f3",
          1212 => x"3d0d7f61",
          1213 => x"63028c05",
          1214 => x"80cf0533",
          1215 => x"73731568",
          1216 => x"415f5c5c",
          1217 => x"5e5e5e7a",
          1218 => x"5281eee8",
          1219 => x"51aecc3f",
          1220 => x"81eef051",
          1221 => x"a8d53f80",
          1222 => x"55747927",
          1223 => x"80f4387b",
          1224 => x"902e8938",
          1225 => x"7ba02ea4",
          1226 => x"3880c139",
          1227 => x"74185372",
          1228 => x"7a278d38",
          1229 => x"72225281",
          1230 => x"eef451ae",
          1231 => x"9e3f8839",
          1232 => x"81ef8051",
          1233 => x"a8a53f82",
          1234 => x"1555bf39",
          1235 => x"74185372",
          1236 => x"7a278d38",
          1237 => x"72085281",
          1238 => x"eee851ad",
          1239 => x"fe3f8839",
          1240 => x"81eefc51",
          1241 => x"a8853f84",
          1242 => x"15559f39",
          1243 => x"74185372",
          1244 => x"7a278d38",
          1245 => x"72335281",
          1246 => x"ef8851ad",
          1247 => x"de3f8839",
          1248 => x"81ef9051",
          1249 => x"a7e53f81",
          1250 => x"1555a051",
          1251 => x"a7803fff",
          1252 => x"883981ef",
          1253 => x"9451a7d3",
          1254 => x"3f805574",
          1255 => x"7927bb38",
          1256 => x"74187033",
          1257 => x"55538056",
          1258 => x"727a2783",
          1259 => x"38815680",
          1260 => x"539f7427",
          1261 => x"83388153",
          1262 => x"75730670",
          1263 => x"81ff0651",
          1264 => x"5372802e",
          1265 => x"8b387380",
          1266 => x"fe268538",
          1267 => x"73518339",
          1268 => x"a051a6ba",
          1269 => x"3f811555",
          1270 => x"c23981ef",
          1271 => x"9851a78b",
          1272 => x"3f781879",
          1273 => x"1c5c589b",
          1274 => x"fb3f8285",
          1275 => x"ec08982b",
          1276 => x"70982c51",
          1277 => x"5776a02e",
          1278 => x"098106ae",
          1279 => x"389be53f",
          1280 => x"8285ec08",
          1281 => x"982b7098",
          1282 => x"2c70a032",
          1283 => x"70098105",
          1284 => x"729b3270",
          1285 => x"09810570",
          1286 => x"72077375",
          1287 => x"07065158",
          1288 => x"58595751",
          1289 => x"57807324",
          1290 => x"d438769b",
          1291 => x"2e098106",
          1292 => x"85388053",
          1293 => x"8c397c1e",
          1294 => x"53727826",
          1295 => x"fdc938ff",
          1296 => x"53728285",
          1297 => x"ec0c8f3d",
          1298 => x"0d04fc3d",
          1299 => x"0d029b05",
          1300 => x"3381ef9c",
          1301 => x"5381efa0",
          1302 => x"5255abff",
          1303 => x"3f8284c4",
          1304 => x"2251a4d1",
          1305 => x"3f81efac",
          1306 => x"5481efb8",
          1307 => x"538284c5",
          1308 => x"335281ef",
          1309 => x"c051abe3",
          1310 => x"3f74802e",
          1311 => x"8438a086",
          1312 => x"3f863d0d",
          1313 => x"04fe3d0d",
          1314 => x"87c09680",
          1315 => x"0853a4ec",
          1316 => x"3f815196",
          1317 => x"eb3f81ef",
          1318 => x"dc5198e0",
          1319 => x"3f805196",
          1320 => x"df3f7281",
          1321 => x"2a708106",
          1322 => x"51527180",
          1323 => x"2e923881",
          1324 => x"5196cd3f",
          1325 => x"81eff451",
          1326 => x"98c23f80",
          1327 => x"5196c13f",
          1328 => x"72822a70",
          1329 => x"81065152",
          1330 => x"71802e92",
          1331 => x"38815196",
          1332 => x"af3f81f0",
          1333 => x"885198a4",
          1334 => x"3f805196",
          1335 => x"a33f7283",
          1336 => x"2a708106",
          1337 => x"51527180",
          1338 => x"2e923881",
          1339 => x"5196913f",
          1340 => x"81f09851",
          1341 => x"98863f80",
          1342 => x"5196853f",
          1343 => x"72842a70",
          1344 => x"81065152",
          1345 => x"71802e92",
          1346 => x"38815195",
          1347 => x"f33f81f0",
          1348 => x"ac5197e8",
          1349 => x"3f805195",
          1350 => x"e73f7285",
          1351 => x"2a708106",
          1352 => x"51527180",
          1353 => x"2e923881",
          1354 => x"5195d53f",
          1355 => x"81f0c051",
          1356 => x"97ca3f80",
          1357 => x"5195c93f",
          1358 => x"72862a70",
          1359 => x"81065152",
          1360 => x"71802e92",
          1361 => x"38815195",
          1362 => x"b73f81f0",
          1363 => x"d45197ac",
          1364 => x"3f805195",
          1365 => x"ab3f7287",
          1366 => x"2a708106",
          1367 => x"51527180",
          1368 => x"2e923881",
          1369 => x"5195993f",
          1370 => x"81f0e851",
          1371 => x"978e3f80",
          1372 => x"51958d3f",
          1373 => x"72882a70",
          1374 => x"81065152",
          1375 => x"71802e92",
          1376 => x"38815194",
          1377 => x"fb3f81f0",
          1378 => x"fc5196f0",
          1379 => x"3f805194",
          1380 => x"ef3fa2f0",
          1381 => x"3f843d0d",
          1382 => x"04fb3d0d",
          1383 => x"77028405",
          1384 => x"a3053370",
          1385 => x"55565680",
          1386 => x"527551ed",
          1387 => x"c03f0b0b",
          1388 => x"8280e833",
          1389 => x"5473ab38",
          1390 => x"815381f1",
          1391 => x"bc52829c",
          1392 => x"cc5180fe",
          1393 => x"f73f8285",
          1394 => x"ec080981",
          1395 => x"05708285",
          1396 => x"ec080780",
          1397 => x"25827131",
          1398 => x"51515473",
          1399 => x"0b0b8280",
          1400 => x"e8340b0b",
          1401 => x"8280e833",
          1402 => x"5473812e",
          1403 => x"098106af",
          1404 => x"38829ccc",
          1405 => x"53745275",
          1406 => x"5181b9c4",
          1407 => x"3f8285ec",
          1408 => x"08802e8b",
          1409 => x"388285ec",
          1410 => x"0851a2df",
          1411 => x"3f913982",
          1412 => x"9ccc5181",
          1413 => x"8b993f82",
          1414 => x"0b0b0b82",
          1415 => x"80e8340b",
          1416 => x"0b8280e8",
          1417 => x"33547382",
          1418 => x"2e098106",
          1419 => x"8c3881f1",
          1420 => x"cc537452",
          1421 => x"7551b592",
          1422 => x"3f800b82",
          1423 => x"85ec0c87",
          1424 => x"3d0d04ce",
          1425 => x"3d0d8070",
          1426 => x"71829cc8",
          1427 => x"0c5f5d81",
          1428 => x"527c5180",
          1429 => x"cd933f82",
          1430 => x"85ec0881",
          1431 => x"ff065978",
          1432 => x"7d2e0981",
          1433 => x"06a13881",
          1434 => x"f1d45296",
          1435 => x"3d705259",
          1436 => x"a7ff3f7c",
          1437 => x"53785282",
          1438 => x"86f85180",
          1439 => x"fcdd3f82",
          1440 => x"85ec087d",
          1441 => x"2e883881",
          1442 => x"f1d8518d",
          1443 => x"8a398170",
          1444 => x"5f5d81f2",
          1445 => x"9051a1d3",
          1446 => x"3f963d70",
          1447 => x"465a80f8",
          1448 => x"527951fd",
          1449 => x"f43fb43d",
          1450 => x"ff840551",
          1451 => x"f3d43f82",
          1452 => x"85ec0890",
          1453 => x"2b70902c",
          1454 => x"51597880",
          1455 => x"c22e879c",
          1456 => x"387880c2",
          1457 => x"24b23878",
          1458 => x"bd2e81d1",
          1459 => x"3878bd24",
          1460 => x"90387880",
          1461 => x"2effbb38",
          1462 => x"78bc2e80",
          1463 => x"da388abb",
          1464 => x"397880c0",
          1465 => x"2e839438",
          1466 => x"7880c024",
          1467 => x"85cd3878",
          1468 => x"bf2e828a",
          1469 => x"388aa439",
          1470 => x"7880f92e",
          1471 => x"89c33878",
          1472 => x"80f92492",
          1473 => x"387880c3",
          1474 => x"2e87fa38",
          1475 => x"7880f82e",
          1476 => x"898c388a",
          1477 => x"86397881",
          1478 => x"832e89ed",
          1479 => x"38788183",
          1480 => x"248b3878",
          1481 => x"81822e89",
          1482 => x"d33889ef",
          1483 => x"39788185",
          1484 => x"2e89e238",
          1485 => x"89e539b4",
          1486 => x"3dff8011",
          1487 => x"53ff8405",
          1488 => x"51a8903f",
          1489 => x"8285ec08",
          1490 => x"802efec6",
          1491 => x"38b43dfe",
          1492 => x"fc1153ff",
          1493 => x"840551a7",
          1494 => x"fa3f8285",
          1495 => x"ec08802e",
          1496 => x"feb038b4",
          1497 => x"3dfef811",
          1498 => x"53ff8405",
          1499 => x"51a7e43f",
          1500 => x"8285ec08",
          1501 => x"86388285",
          1502 => x"ec084281",
          1503 => x"f294519f",
          1504 => x"ea3f6363",
          1505 => x"5c5a797b",
          1506 => x"2781e938",
          1507 => x"6159787a",
          1508 => x"7084055c",
          1509 => x"0c7a7a26",
          1510 => x"f53881d8",
          1511 => x"39b43dff",
          1512 => x"801153ff",
          1513 => x"840551a7",
          1514 => x"aa3f8285",
          1515 => x"ec08802e",
          1516 => x"fde038b4",
          1517 => x"3dfefc11",
          1518 => x"53ff8405",
          1519 => x"51a7943f",
          1520 => x"8285ec08",
          1521 => x"802efdca",
          1522 => x"38b43dfe",
          1523 => x"f81153ff",
          1524 => x"840551a6",
          1525 => x"fe3f8285",
          1526 => x"ec08802e",
          1527 => x"fdb43881",
          1528 => x"f2a4519f",
          1529 => x"863f635a",
          1530 => x"79632781",
          1531 => x"87386159",
          1532 => x"79708105",
          1533 => x"5b337934",
          1534 => x"61810542",
          1535 => x"eb39b43d",
          1536 => x"ff801153",
          1537 => x"ff840551",
          1538 => x"a6c93f82",
          1539 => x"85ec0880",
          1540 => x"2efcff38",
          1541 => x"b43dfefc",
          1542 => x"1153ff84",
          1543 => x"0551a6b3",
          1544 => x"3f8285ec",
          1545 => x"08802efc",
          1546 => x"e938b43d",
          1547 => x"fef81153",
          1548 => x"ff840551",
          1549 => x"a69d3f82",
          1550 => x"85ec0880",
          1551 => x"2efcd338",
          1552 => x"81f2b051",
          1553 => x"9ea53f63",
          1554 => x"5a796327",
          1555 => x"a7386170",
          1556 => x"337b335e",
          1557 => x"5a5b787c",
          1558 => x"2e913878",
          1559 => x"557a5479",
          1560 => x"33537952",
          1561 => x"81f2c051",
          1562 => x"a3f13f81",
          1563 => x"1a628105",
          1564 => x"435ad639",
          1565 => x"81f2d851",
          1566 => x"82bb39b4",
          1567 => x"3dff8011",
          1568 => x"53ff8405",
          1569 => x"51a5cc3f",
          1570 => x"8285ec08",
          1571 => x"80df3882",
          1572 => x"84d83359",
          1573 => x"78802e89",
          1574 => x"38828490",
          1575 => x"084480cd",
          1576 => x"398284d9",
          1577 => x"33597880",
          1578 => x"2e883882",
          1579 => x"84980844",
          1580 => x"bc398284",
          1581 => x"da335978",
          1582 => x"802e8838",
          1583 => x"8284a008",
          1584 => x"44ab3982",
          1585 => x"84db3359",
          1586 => x"78802e88",
          1587 => x"388284a8",
          1588 => x"08449a39",
          1589 => x"8284d633",
          1590 => x"5978802e",
          1591 => x"88388284",
          1592 => x"b0084489",
          1593 => x"398284c0",
          1594 => x"08fc8005",
          1595 => x"44b43dfe",
          1596 => x"fc1153ff",
          1597 => x"840551a4",
          1598 => x"da3f8285",
          1599 => x"ec0880de",
          1600 => x"388284d8",
          1601 => x"33597880",
          1602 => x"2e893882",
          1603 => x"84940843",
          1604 => x"80cc3982",
          1605 => x"84d93359",
          1606 => x"78802e88",
          1607 => x"3882849c",
          1608 => x"0843bb39",
          1609 => x"8284da33",
          1610 => x"5978802e",
          1611 => x"88388284",
          1612 => x"a40843aa",
          1613 => x"398284db",
          1614 => x"33597880",
          1615 => x"2e883882",
          1616 => x"84ac0843",
          1617 => x"99398284",
          1618 => x"d6335978",
          1619 => x"802e8838",
          1620 => x"8284b408",
          1621 => x"43883982",
          1622 => x"84c00888",
          1623 => x"0543b43d",
          1624 => x"fef81153",
          1625 => x"ff840551",
          1626 => x"a3e93f82",
          1627 => x"85ec0880",
          1628 => x"2ea93880",
          1629 => x"625c5c7a",
          1630 => x"882e8338",
          1631 => x"815c7a90",
          1632 => x"32700981",
          1633 => x"05707207",
          1634 => x"9f2a707f",
          1635 => x"0651515a",
          1636 => x"5a78802e",
          1637 => x"88387aa0",
          1638 => x"2e833888",
          1639 => x"4281f2dc",
          1640 => x"519bc83f",
          1641 => x"a0556354",
          1642 => x"61536252",
          1643 => x"6351f2bf",
          1644 => x"3f81f2ec",
          1645 => x"519bb43f",
          1646 => x"f9d839b4",
          1647 => x"3dff8011",
          1648 => x"53ff8405",
          1649 => x"51a38c3f",
          1650 => x"8285ec08",
          1651 => x"802ef9c2",
          1652 => x"38b43dfe",
          1653 => x"fc1153ff",
          1654 => x"840551a2",
          1655 => x"f63f8285",
          1656 => x"ec08802e",
          1657 => x"a4386359",
          1658 => x"0280cb05",
          1659 => x"33793463",
          1660 => x"810544b4",
          1661 => x"3dfefc11",
          1662 => x"53ff8405",
          1663 => x"51a2d43f",
          1664 => x"8285ec08",
          1665 => x"e138f98a",
          1666 => x"39637033",
          1667 => x"545281f2",
          1668 => x"f851a0c7",
          1669 => x"3f80f852",
          1670 => x"7951a199",
          1671 => x"3f794579",
          1672 => x"335978ae",
          1673 => x"2ef8eb38",
          1674 => x"9f79279f",
          1675 => x"38b43dfe",
          1676 => x"fc1153ff",
          1677 => x"840551a2",
          1678 => x"9a3f8285",
          1679 => x"ec08802e",
          1680 => x"91386359",
          1681 => x"0280cb05",
          1682 => x"33793463",
          1683 => x"810544ff",
          1684 => x"b83981f3",
          1685 => x"84519a93",
          1686 => x"3fffae39",
          1687 => x"b43dfef4",
          1688 => x"1153ff84",
          1689 => x"0551a3e7",
          1690 => x"3f8285ec",
          1691 => x"08802ef8",
          1692 => x"a138b43d",
          1693 => x"fef01153",
          1694 => x"ff840551",
          1695 => x"a3d13f82",
          1696 => x"85ec0880",
          1697 => x"2ea53860",
          1698 => x"5902be05",
          1699 => x"22797082",
          1700 => x"055b2378",
          1701 => x"41b43dfe",
          1702 => x"f01153ff",
          1703 => x"840551a3",
          1704 => x"ae3f8285",
          1705 => x"ec08e038",
          1706 => x"f7e83960",
          1707 => x"70225452",
          1708 => x"81f38c51",
          1709 => x"9fa53f80",
          1710 => x"f8527951",
          1711 => x"9ff73f79",
          1712 => x"45793359",
          1713 => x"78ae2ef7",
          1714 => x"c938789f",
          1715 => x"26873860",
          1716 => x"820541d7",
          1717 => x"39b43dfe",
          1718 => x"f01153ff",
          1719 => x"840551a2",
          1720 => x"ee3f8285",
          1721 => x"ec08802e",
          1722 => x"92386059",
          1723 => x"02be0522",
          1724 => x"79708205",
          1725 => x"5b237841",
          1726 => x"ffb13981",
          1727 => x"f3845198",
          1728 => x"ea3fffa7",
          1729 => x"39b43dfe",
          1730 => x"f41153ff",
          1731 => x"840551a2",
          1732 => x"be3f8285",
          1733 => x"ec08802e",
          1734 => x"f6f838b4",
          1735 => x"3dfef011",
          1736 => x"53ff8405",
          1737 => x"51a2a83f",
          1738 => x"8285ec08",
          1739 => x"802ea038",
          1740 => x"6060710c",
          1741 => x"59608405",
          1742 => x"41b43dfe",
          1743 => x"f01153ff",
          1744 => x"840551a2",
          1745 => x"8a3f8285",
          1746 => x"ec08e538",
          1747 => x"f6c43960",
          1748 => x"70085452",
          1749 => x"81f39851",
          1750 => x"9e813f80",
          1751 => x"f8527951",
          1752 => x"9ed33f79",
          1753 => x"45793359",
          1754 => x"78ae2ef6",
          1755 => x"a5389f79",
          1756 => x"279b38b4",
          1757 => x"3dfef011",
          1758 => x"53ff8405",
          1759 => x"51a1d03f",
          1760 => x"8285ec08",
          1761 => x"802e8d38",
          1762 => x"6060710c",
          1763 => x"59608405",
          1764 => x"41ffbc39",
          1765 => x"81f38451",
          1766 => x"97d13fff",
          1767 => x"b239b43d",
          1768 => x"ff801153",
          1769 => x"ff840551",
          1770 => x"9fa93f82",
          1771 => x"85ec0880",
          1772 => x"2ef5df38",
          1773 => x"635281f3",
          1774 => x"a4519d9f",
          1775 => x"3f635978",
          1776 => x"04b43dff",
          1777 => x"801153ff",
          1778 => x"8405519f",
          1779 => x"863f8285",
          1780 => x"ec08802e",
          1781 => x"f5bc3863",
          1782 => x"5281f3c0",
          1783 => x"519cfc3f",
          1784 => x"6359782d",
          1785 => x"8285ec08",
          1786 => x"802ef5a6",
          1787 => x"388285ec",
          1788 => x"085281f3",
          1789 => x"dc519ce3",
          1790 => x"3ff59739",
          1791 => x"81f3f851",
          1792 => x"96e93fdb",
          1793 => x"963ff58a",
          1794 => x"3981f494",
          1795 => x"5196dc3f",
          1796 => x"8059ffab",
          1797 => x"3990ef3f",
          1798 => x"f4f83979",
          1799 => x"45793359",
          1800 => x"78802ef4",
          1801 => x"ed387d7d",
          1802 => x"06597880",
          1803 => x"2e81d038",
          1804 => x"b43dff84",
          1805 => x"055183b5",
          1806 => x"3f8285ec",
          1807 => x"085c815b",
          1808 => x"7a822eb1",
          1809 => x"387a8224",
          1810 => x"89387a81",
          1811 => x"2e8c3880",
          1812 => x"ca397a83",
          1813 => x"2eae3880",
          1814 => x"c23981f4",
          1815 => x"a8567b55",
          1816 => x"81f4ac54",
          1817 => x"805381f4",
          1818 => x"b052b43d",
          1819 => x"ffb00551",
          1820 => x"9bff3fb8",
          1821 => x"3981f4d0",
          1822 => x"52b43dff",
          1823 => x"b005519b",
          1824 => x"f03fa939",
          1825 => x"7b5581f4",
          1826 => x"ac548053",
          1827 => x"81f4c052",
          1828 => x"b43dffb0",
          1829 => x"05519bd9",
          1830 => x"3f92397b",
          1831 => x"54805381",
          1832 => x"f4cc52b4",
          1833 => x"3dffb005",
          1834 => x"519bc63f",
          1835 => x"82849058",
          1836 => x"8285fc57",
          1837 => x"80566455",
          1838 => x"805482a0",
          1839 => x"805382a0",
          1840 => x"8052b43d",
          1841 => x"ffb00551",
          1842 => x"ebdc3f82",
          1843 => x"85ec0882",
          1844 => x"85ec0809",
          1845 => x"70098105",
          1846 => x"70720780",
          1847 => x"25515b5b",
          1848 => x"5f805a7a",
          1849 => x"83268338",
          1850 => x"815a787a",
          1851 => x"06597880",
          1852 => x"2e8d3881",
          1853 => x"1b7081ff",
          1854 => x"065c597a",
          1855 => x"fec2387d",
          1856 => x"81327d81",
          1857 => x"32075978",
          1858 => x"8a387eff",
          1859 => x"2e098106",
          1860 => x"f3803881",
          1861 => x"f4d4519a",
          1862 => x"c23ff2f6",
          1863 => x"39fc3d0d",
          1864 => x"800b8285",
          1865 => x"fc3487c0",
          1866 => x"948c7008",
          1867 => x"54558784",
          1868 => x"80527251",
          1869 => x"e3d43f82",
          1870 => x"85ec0890",
          1871 => x"2b750855",
          1872 => x"53878480",
          1873 => x"527351e3",
          1874 => x"c13f7282",
          1875 => x"85ec0807",
          1876 => x"750c87c0",
          1877 => x"949c7008",
          1878 => x"54558784",
          1879 => x"80527251",
          1880 => x"e3a83f82",
          1881 => x"85ec0890",
          1882 => x"2b750855",
          1883 => x"53878480",
          1884 => x"527351e3",
          1885 => x"953f7282",
          1886 => x"85ec0807",
          1887 => x"750c8c80",
          1888 => x"830b87c0",
          1889 => x"94840c8c",
          1890 => x"80830b87",
          1891 => x"c094940c",
          1892 => x"80c09a0b",
          1893 => x"829cf40c",
          1894 => x"80c3950b",
          1895 => x"829cf80c",
          1896 => x"89983f92",
          1897 => x"d73f81f4",
          1898 => x"e45193bf",
          1899 => x"3f81f4f0",
          1900 => x"5193b83f",
          1901 => x"a9855192",
          1902 => x"be3f8151",
          1903 => x"ed8c3ff1",
          1904 => x"823f8004",
          1905 => x"fe3d0d80",
          1906 => x"52835371",
          1907 => x"882b5287",
          1908 => x"c43f8285",
          1909 => x"ec0881ff",
          1910 => x"067207ff",
          1911 => x"14545272",
          1912 => x"8025e838",
          1913 => x"718285ec",
          1914 => x"0c843d0d",
          1915 => x"04fc3d0d",
          1916 => x"76700854",
          1917 => x"55807352",
          1918 => x"5472742e",
          1919 => x"818c3872",
          1920 => x"335170a0",
          1921 => x"2e098106",
          1922 => x"86388113",
          1923 => x"53f13972",
          1924 => x"335170a2",
          1925 => x"2e098106",
          1926 => x"86388113",
          1927 => x"53815472",
          1928 => x"5273812e",
          1929 => x"0981069f",
          1930 => x"38843981",
          1931 => x"12528072",
          1932 => x"33525470",
          1933 => x"a22e8338",
          1934 => x"81547080",
          1935 => x"2e9d3873",
          1936 => x"ea389839",
          1937 => x"81125280",
          1938 => x"72335254",
          1939 => x"70a02e83",
          1940 => x"38815470",
          1941 => x"802e8438",
          1942 => x"73ea3880",
          1943 => x"72335254",
          1944 => x"70a02e09",
          1945 => x"81068338",
          1946 => x"815470a2",
          1947 => x"32700981",
          1948 => x"05708025",
          1949 => x"76075151",
          1950 => x"5170802e",
          1951 => x"88388072",
          1952 => x"70810554",
          1953 => x"3471750c",
          1954 => x"72517082",
          1955 => x"85ec0c86",
          1956 => x"3d0d04fc",
          1957 => x"3d0d7653",
          1958 => x"7208802e",
          1959 => x"9138863d",
          1960 => x"fc055272",
          1961 => x"519ba83f",
          1962 => x"8285ec08",
          1963 => x"85388053",
          1964 => x"83397453",
          1965 => x"728285ec",
          1966 => x"0c863d0d",
          1967 => x"04fc3d0d",
          1968 => x"76821133",
          1969 => x"ff055253",
          1970 => x"8152708b",
          1971 => x"26819838",
          1972 => x"831333ff",
          1973 => x"05518252",
          1974 => x"709e2681",
          1975 => x"8a388413",
          1976 => x"33518352",
          1977 => x"70972680",
          1978 => x"fe388513",
          1979 => x"33518452",
          1980 => x"70bb2680",
          1981 => x"f2388613",
          1982 => x"33518552",
          1983 => x"70bb2680",
          1984 => x"e6388813",
          1985 => x"22558652",
          1986 => x"7487e726",
          1987 => x"80d9388a",
          1988 => x"13225487",
          1989 => x"527387e7",
          1990 => x"2680cc38",
          1991 => x"810b87c0",
          1992 => x"989c0c72",
          1993 => x"2287c098",
          1994 => x"bc0c8213",
          1995 => x"3387c098",
          1996 => x"b80c8313",
          1997 => x"3387c098",
          1998 => x"b40c8413",
          1999 => x"3387c098",
          2000 => x"b00c8513",
          2001 => x"3387c098",
          2002 => x"ac0c8613",
          2003 => x"3387c098",
          2004 => x"a80c7487",
          2005 => x"c098a40c",
          2006 => x"7387c098",
          2007 => x"a00c800b",
          2008 => x"87c0989c",
          2009 => x"0c805271",
          2010 => x"8285ec0c",
          2011 => x"863d0d04",
          2012 => x"f33d0d7f",
          2013 => x"5b87c098",
          2014 => x"9c5d817d",
          2015 => x"0c87c098",
          2016 => x"bc085e7d",
          2017 => x"7b2387c0",
          2018 => x"98b8085a",
          2019 => x"79821c34",
          2020 => x"87c098b4",
          2021 => x"085a7983",
          2022 => x"1c3487c0",
          2023 => x"98b0085a",
          2024 => x"79841c34",
          2025 => x"87c098ac",
          2026 => x"085a7985",
          2027 => x"1c3487c0",
          2028 => x"98a8085a",
          2029 => x"79861c34",
          2030 => x"87c098a4",
          2031 => x"085c7b88",
          2032 => x"1c2387c0",
          2033 => x"98a0085a",
          2034 => x"798a1c23",
          2035 => x"807d0c79",
          2036 => x"83ffff06",
          2037 => x"597b83ff",
          2038 => x"ff065886",
          2039 => x"1b335785",
          2040 => x"1b335684",
          2041 => x"1b335583",
          2042 => x"1b335482",
          2043 => x"1b33537d",
          2044 => x"83ffff06",
          2045 => x"5281f588",
          2046 => x"5194e03f",
          2047 => x"8f3d0d04",
          2048 => x"ff3d0d02",
          2049 => x"8f053370",
          2050 => x"09810570",
          2051 => x"9f2a5152",
          2052 => x"52708284",
          2053 => x"8c34833d",
          2054 => x"0d04fb3d",
          2055 => x"0d778284",
          2056 => x"8c337081",
          2057 => x"ff065755",
          2058 => x"5687c094",
          2059 => x"84517480",
          2060 => x"2e863887",
          2061 => x"c0949451",
          2062 => x"70087096",
          2063 => x"2a708106",
          2064 => x"53545270",
          2065 => x"802e8c38",
          2066 => x"71912a70",
          2067 => x"81065151",
          2068 => x"70d73872",
          2069 => x"81327081",
          2070 => x"06515170",
          2071 => x"802e8d38",
          2072 => x"71932a70",
          2073 => x"81065151",
          2074 => x"70ffbe38",
          2075 => x"7381ff06",
          2076 => x"5187c094",
          2077 => x"80527080",
          2078 => x"2e863887",
          2079 => x"c0949052",
          2080 => x"75720c75",
          2081 => x"8285ec0c",
          2082 => x"873d0d04",
          2083 => x"fb3d0d02",
          2084 => x"9f053382",
          2085 => x"848c3370",
          2086 => x"81ff0657",
          2087 => x"555687c0",
          2088 => x"94845174",
          2089 => x"802e8638",
          2090 => x"87c09494",
          2091 => x"51700870",
          2092 => x"962a7081",
          2093 => x"06535452",
          2094 => x"70802e8c",
          2095 => x"3871912a",
          2096 => x"70810651",
          2097 => x"5170d738",
          2098 => x"72813270",
          2099 => x"81065151",
          2100 => x"70802e8d",
          2101 => x"3871932a",
          2102 => x"70810651",
          2103 => x"5170ffbe",
          2104 => x"387381ff",
          2105 => x"065187c0",
          2106 => x"94805270",
          2107 => x"802e8638",
          2108 => x"87c09490",
          2109 => x"5275720c",
          2110 => x"873d0d04",
          2111 => x"f93d0d79",
          2112 => x"54807433",
          2113 => x"7081ff06",
          2114 => x"53535770",
          2115 => x"772e80fc",
          2116 => x"387181ff",
          2117 => x"06811582",
          2118 => x"848c3370",
          2119 => x"81ff0659",
          2120 => x"57555887",
          2121 => x"c0948451",
          2122 => x"75802e86",
          2123 => x"3887c094",
          2124 => x"94517008",
          2125 => x"70962a70",
          2126 => x"81065354",
          2127 => x"5270802e",
          2128 => x"8c387191",
          2129 => x"2a708106",
          2130 => x"515170d7",
          2131 => x"38728132",
          2132 => x"70810651",
          2133 => x"5170802e",
          2134 => x"8d387193",
          2135 => x"2a708106",
          2136 => x"515170ff",
          2137 => x"be387481",
          2138 => x"ff065187",
          2139 => x"c0948052",
          2140 => x"70802e86",
          2141 => x"3887c094",
          2142 => x"90527772",
          2143 => x"0c811774",
          2144 => x"337081ff",
          2145 => x"06535357",
          2146 => x"70ff8638",
          2147 => x"768285ec",
          2148 => x"0c893d0d",
          2149 => x"04fe3d0d",
          2150 => x"82848c33",
          2151 => x"7081ff06",
          2152 => x"545287c0",
          2153 => x"94845172",
          2154 => x"802e8638",
          2155 => x"87c09494",
          2156 => x"51700870",
          2157 => x"822a7081",
          2158 => x"06515151",
          2159 => x"70802ee2",
          2160 => x"387181ff",
          2161 => x"065187c0",
          2162 => x"94805270",
          2163 => x"802e8638",
          2164 => x"87c09490",
          2165 => x"52710870",
          2166 => x"81ff0682",
          2167 => x"85ec0c51",
          2168 => x"843d0d04",
          2169 => x"fe3d0d82",
          2170 => x"848c3370",
          2171 => x"81ff0652",
          2172 => x"5387c094",
          2173 => x"84527080",
          2174 => x"2e863887",
          2175 => x"c0949452",
          2176 => x"71087082",
          2177 => x"2a708106",
          2178 => x"515151ff",
          2179 => x"5270802e",
          2180 => x"a0387281",
          2181 => x"ff065187",
          2182 => x"c0948052",
          2183 => x"70802e86",
          2184 => x"3887c094",
          2185 => x"90527108",
          2186 => x"70982b70",
          2187 => x"982c5153",
          2188 => x"51718285",
          2189 => x"ec0c843d",
          2190 => x"0d04ff3d",
          2191 => x"0d87c09e",
          2192 => x"8008709c",
          2193 => x"2a8a0651",
          2194 => x"5170802e",
          2195 => x"84b43887",
          2196 => x"c09ea408",
          2197 => x"8284900c",
          2198 => x"87c09ea8",
          2199 => x"08828494",
          2200 => x"0c87c09e",
          2201 => x"94088284",
          2202 => x"980c87c0",
          2203 => x"9e980882",
          2204 => x"849c0c87",
          2205 => x"c09e9c08",
          2206 => x"8284a00c",
          2207 => x"87c09ea0",
          2208 => x"088284a4",
          2209 => x"0c87c09e",
          2210 => x"ac088284",
          2211 => x"a80c87c0",
          2212 => x"9eb00882",
          2213 => x"84ac0c87",
          2214 => x"c09eb408",
          2215 => x"8284b00c",
          2216 => x"87c09eb8",
          2217 => x"088284b4",
          2218 => x"0c87c09e",
          2219 => x"bc088284",
          2220 => x"b80c87c0",
          2221 => x"9ec00882",
          2222 => x"84bc0c87",
          2223 => x"c09ec408",
          2224 => x"8284c00c",
          2225 => x"87c09e80",
          2226 => x"08517082",
          2227 => x"84c42387",
          2228 => x"c09e8408",
          2229 => x"8284c80c",
          2230 => x"87c09e88",
          2231 => x"088284cc",
          2232 => x"0c87c09e",
          2233 => x"8c088284",
          2234 => x"d00c810b",
          2235 => x"8284d434",
          2236 => x"800b87c0",
          2237 => x"9e900870",
          2238 => x"84800a06",
          2239 => x"51525270",
          2240 => x"802e8338",
          2241 => x"81527182",
          2242 => x"84d53480",
          2243 => x"0b87c09e",
          2244 => x"90087088",
          2245 => x"800a0651",
          2246 => x"52527080",
          2247 => x"2e833881",
          2248 => x"52718284",
          2249 => x"d634800b",
          2250 => x"87c09e90",
          2251 => x"08709080",
          2252 => x"0a065152",
          2253 => x"5270802e",
          2254 => x"83388152",
          2255 => x"718284d7",
          2256 => x"34800b87",
          2257 => x"c09e9008",
          2258 => x"70888080",
          2259 => x"06515252",
          2260 => x"70802e83",
          2261 => x"38815271",
          2262 => x"8284d834",
          2263 => x"800b87c0",
          2264 => x"9e900870",
          2265 => x"a0808006",
          2266 => x"51525270",
          2267 => x"802e8338",
          2268 => x"81527182",
          2269 => x"84d93480",
          2270 => x"0b87c09e",
          2271 => x"90087090",
          2272 => x"80800651",
          2273 => x"52527080",
          2274 => x"2e833881",
          2275 => x"52718284",
          2276 => x"da34800b",
          2277 => x"87c09e90",
          2278 => x"08708480",
          2279 => x"80065152",
          2280 => x"5270802e",
          2281 => x"83388152",
          2282 => x"718284db",
          2283 => x"34800b87",
          2284 => x"c09e9008",
          2285 => x"70828080",
          2286 => x"06515252",
          2287 => x"70802e83",
          2288 => x"38815271",
          2289 => x"8284dc34",
          2290 => x"800b87c0",
          2291 => x"9e900870",
          2292 => x"81808006",
          2293 => x"51525270",
          2294 => x"802e8338",
          2295 => x"81527182",
          2296 => x"84dd3480",
          2297 => x"0b87c09e",
          2298 => x"90087080",
          2299 => x"c0800651",
          2300 => x"52527080",
          2301 => x"2e833881",
          2302 => x"52718284",
          2303 => x"de34800b",
          2304 => x"87c09e90",
          2305 => x"0870a080",
          2306 => x"06515252",
          2307 => x"70802e83",
          2308 => x"38815271",
          2309 => x"8284df34",
          2310 => x"87c09e90",
          2311 => x"08709880",
          2312 => x"06708a2a",
          2313 => x"51515170",
          2314 => x"8284e034",
          2315 => x"800b87c0",
          2316 => x"9e900870",
          2317 => x"84800651",
          2318 => x"52527080",
          2319 => x"2e833881",
          2320 => x"52718284",
          2321 => x"e13487c0",
          2322 => x"9e900870",
          2323 => x"83f00670",
          2324 => x"842a5151",
          2325 => x"51708284",
          2326 => x"e234800b",
          2327 => x"87c09e90",
          2328 => x"08708806",
          2329 => x"51525270",
          2330 => x"802e8338",
          2331 => x"81527182",
          2332 => x"84e33487",
          2333 => x"c09e9008",
          2334 => x"70870651",
          2335 => x"51708284",
          2336 => x"e434833d",
          2337 => x"0d04fc3d",
          2338 => x"0d81f5a0",
          2339 => x"5185dc3f",
          2340 => x"8284d433",
          2341 => x"5473802e",
          2342 => x"883881f5",
          2343 => x"b45185cb",
          2344 => x"3f81f5c8",
          2345 => x"5185c43f",
          2346 => x"8284d633",
          2347 => x"5473802e",
          2348 => x"93388284",
          2349 => x"b0088284",
          2350 => x"b4081154",
          2351 => x"5281f5e0",
          2352 => x"518b983f",
          2353 => x"8284db33",
          2354 => x"5473802e",
          2355 => x"93388284",
          2356 => x"a8088284",
          2357 => x"ac081154",
          2358 => x"5281f5fc",
          2359 => x"518afc3f",
          2360 => x"8284d833",
          2361 => x"5473802e",
          2362 => x"93388284",
          2363 => x"90088284",
          2364 => x"94081154",
          2365 => x"5281f698",
          2366 => x"518ae03f",
          2367 => x"8284d933",
          2368 => x"5473802e",
          2369 => x"93388284",
          2370 => x"98088284",
          2371 => x"9c081154",
          2372 => x"5281f6b4",
          2373 => x"518ac43f",
          2374 => x"8284da33",
          2375 => x"5473802e",
          2376 => x"93388284",
          2377 => x"a0088284",
          2378 => x"a4081154",
          2379 => x"5281f6d0",
          2380 => x"518aa83f",
          2381 => x"8284df33",
          2382 => x"5473802e",
          2383 => x"8d388284",
          2384 => x"e0335281",
          2385 => x"f6ec518a",
          2386 => x"923f8284",
          2387 => x"e3335473",
          2388 => x"802e8d38",
          2389 => x"8284e433",
          2390 => x"5281f78c",
          2391 => x"5189fc3f",
          2392 => x"8284e133",
          2393 => x"5473802e",
          2394 => x"8d388284",
          2395 => x"e2335281",
          2396 => x"f7ac5189",
          2397 => x"e63f8284",
          2398 => x"d5335473",
          2399 => x"802e8838",
          2400 => x"81f7cc51",
          2401 => x"83e53f82",
          2402 => x"84d73354",
          2403 => x"73802e88",
          2404 => x"3881f7e0",
          2405 => x"5183d43f",
          2406 => x"8284dc33",
          2407 => x"5473802e",
          2408 => x"883881f7",
          2409 => x"ec5183c3",
          2410 => x"3f8284dd",
          2411 => x"33547380",
          2412 => x"2e883881",
          2413 => x"f7f85183",
          2414 => x"b23f8284",
          2415 => x"de335473",
          2416 => x"802e8838",
          2417 => x"81f88451",
          2418 => x"83a13f81",
          2419 => x"f8905183",
          2420 => x"9a3f8284",
          2421 => x"b8085281",
          2422 => x"f89c5188",
          2423 => x"fe3f8284",
          2424 => x"bc085281",
          2425 => x"f8c45188",
          2426 => x"f23f8284",
          2427 => x"c0085281",
          2428 => x"f8ec5188",
          2429 => x"e63f81f9",
          2430 => x"945182ef",
          2431 => x"3f8284c4",
          2432 => x"225281f9",
          2433 => x"9c5188d3",
          2434 => x"3f8284c8",
          2435 => x"0855bd84",
          2436 => x"c0527451",
          2437 => x"d1f43f82",
          2438 => x"85ec0854",
          2439 => x"bd84c052",
          2440 => x"8285ec08",
          2441 => x"51d0e33f",
          2442 => x"748285ec",
          2443 => x"08315373",
          2444 => x"5281f9c4",
          2445 => x"5188a43f",
          2446 => x"8284db33",
          2447 => x"5473802e",
          2448 => x"b0388284",
          2449 => x"cc0855bd",
          2450 => x"84c05274",
          2451 => x"51d1bb3f",
          2452 => x"8285ec08",
          2453 => x"54bd84c0",
          2454 => x"528285ec",
          2455 => x"0851d0aa",
          2456 => x"3f748285",
          2457 => x"ec083153",
          2458 => x"735281f9",
          2459 => x"f05187eb",
          2460 => x"3f8284d6",
          2461 => x"33547380",
          2462 => x"2eb03882",
          2463 => x"84d00855",
          2464 => x"bd84c052",
          2465 => x"7451d182",
          2466 => x"3f8285ec",
          2467 => x"0854bd84",
          2468 => x"c0528285",
          2469 => x"ec0851cf",
          2470 => x"f13f7482",
          2471 => x"85ec0831",
          2472 => x"53735281",
          2473 => x"fa9c5187",
          2474 => x"b23f81f2",
          2475 => x"d85181bb",
          2476 => x"3f863d0d",
          2477 => x"04fe3d0d",
          2478 => x"02920533",
          2479 => x"ff055271",
          2480 => x"8426a938",
          2481 => x"71822b52",
          2482 => x"81e8dc12",
          2483 => x"080481fa",
          2484 => x"c8519d39",
          2485 => x"81fad051",
          2486 => x"973981fa",
          2487 => x"d8519139",
          2488 => x"81fae051",
          2489 => x"8b3981fa",
          2490 => x"e4518539",
          2491 => x"81faec51",
          2492 => x"80f93f84",
          2493 => x"3d0d0471",
          2494 => x"88800c04",
          2495 => x"800b87c0",
          2496 => x"96840c04",
          2497 => x"8284e808",
          2498 => x"87c09684",
          2499 => x"0c04fe3d",
          2500 => x"0d029305",
          2501 => x"3353728a",
          2502 => x"2e098106",
          2503 => x"85388d51",
          2504 => x"ed3f829c",
          2505 => x"fc085271",
          2506 => x"802e9038",
          2507 => x"72723482",
          2508 => x"9cfc0881",
          2509 => x"05829cfc",
          2510 => x"0c8f3982",
          2511 => x"9cf40852",
          2512 => x"71802e85",
          2513 => x"38725171",
          2514 => x"2d843d0d",
          2515 => x"04fe3d0d",
          2516 => x"02970533",
          2517 => x"829cf408",
          2518 => x"76829cf4",
          2519 => x"0c5451ff",
          2520 => x"ad3f7282",
          2521 => x"9cf40c84",
          2522 => x"3d0d04fd",
          2523 => x"3d0d7554",
          2524 => x"73337081",
          2525 => x"ff065353",
          2526 => x"71802e8e",
          2527 => x"387281ff",
          2528 => x"06518114",
          2529 => x"54ff873f",
          2530 => x"e739853d",
          2531 => x"0d04fc3d",
          2532 => x"0d77829c",
          2533 => x"f4087882",
          2534 => x"9cf40c56",
          2535 => x"54733370",
          2536 => x"81ff0653",
          2537 => x"5371802e",
          2538 => x"8e387281",
          2539 => x"ff065181",
          2540 => x"1454feda",
          2541 => x"3fe73974",
          2542 => x"829cf40c",
          2543 => x"863d0d04",
          2544 => x"ec3d0d66",
          2545 => x"68595978",
          2546 => x"7081055a",
          2547 => x"33567580",
          2548 => x"2e858438",
          2549 => x"75a52e09",
          2550 => x"810682e4",
          2551 => x"3880707a",
          2552 => x"7081055c",
          2553 => x"33585b5b",
          2554 => x"75b02e09",
          2555 => x"81068538",
          2556 => x"815a8b39",
          2557 => x"75ad2e09",
          2558 => x"81068a38",
          2559 => x"825a7870",
          2560 => x"81055a33",
          2561 => x"5675aa2e",
          2562 => x"09810692",
          2563 => x"38778419",
          2564 => x"71087b70",
          2565 => x"81055d33",
          2566 => x"595d5953",
          2567 => x"9f39d016",
          2568 => x"53728926",
          2569 => x"97387a83",
          2570 => x"2b7b117c",
          2571 => x"1118d005",
          2572 => x"7b708105",
          2573 => x"5d33595d",
          2574 => x"5153e339",
          2575 => x"7580ec32",
          2576 => x"70098105",
          2577 => x"70720780",
          2578 => x"257880cc",
          2579 => x"32700981",
          2580 => x"05707207",
          2581 => x"80257307",
          2582 => x"53545851",
          2583 => x"55537380",
          2584 => x"2e8c3879",
          2585 => x"84077970",
          2586 => x"81055b33",
          2587 => x"575a7580",
          2588 => x"2e83e438",
          2589 => x"755480e0",
          2590 => x"76278938",
          2591 => x"e0167081",
          2592 => x"ff065553",
          2593 => x"7380cf2e",
          2594 => x"81aa3873",
          2595 => x"80cf24a2",
          2596 => x"387380c3",
          2597 => x"2e818e38",
          2598 => x"7380c324",
          2599 => x"8b387380",
          2600 => x"c22e818c",
          2601 => x"38819939",
          2602 => x"7380c42e",
          2603 => x"818a3881",
          2604 => x"8f397380",
          2605 => x"d52e8180",
          2606 => x"387380d5",
          2607 => x"248a3873",
          2608 => x"80d32e8e",
          2609 => x"3880f939",
          2610 => x"7380d82e",
          2611 => x"80ee3880",
          2612 => x"ef397784",
          2613 => x"19710856",
          2614 => x"59538074",
          2615 => x"33545572",
          2616 => x"752e8d38",
          2617 => x"81157015",
          2618 => x"70335154",
          2619 => x"5572f538",
          2620 => x"79812a56",
          2621 => x"90397481",
          2622 => x"16565372",
          2623 => x"7b278f38",
          2624 => x"a051fc8a",
          2625 => x"3f758106",
          2626 => x"5372802e",
          2627 => x"e9387351",
          2628 => x"fcd93f74",
          2629 => x"81165653",
          2630 => x"727b27fd",
          2631 => x"aa38a051",
          2632 => x"fbec3fef",
          2633 => x"39778419",
          2634 => x"83123353",
          2635 => x"59539339",
          2636 => x"825c9539",
          2637 => x"885c9139",
          2638 => x"8a5c8d39",
          2639 => x"905c8939",
          2640 => x"7551fbca",
          2641 => x"3ffd8039",
          2642 => x"79822a70",
          2643 => x"81065153",
          2644 => x"72802e88",
          2645 => x"38778419",
          2646 => x"59538639",
          2647 => x"84187854",
          2648 => x"58720874",
          2649 => x"80c43270",
          2650 => x"09810570",
          2651 => x"72078025",
          2652 => x"51555555",
          2653 => x"7480258f",
          2654 => x"3872802e",
          2655 => x"8a387409",
          2656 => x"81057a90",
          2657 => x"075b5580",
          2658 => x"0b8f3d5e",
          2659 => x"577b5274",
          2660 => x"51cbaa3f",
          2661 => x"8285ec08",
          2662 => x"81ff067c",
          2663 => x"53755254",
          2664 => x"cae83f82",
          2665 => x"85ec0855",
          2666 => x"89742792",
          2667 => x"38a71453",
          2668 => x"7580f82e",
          2669 => x"84388714",
          2670 => x"537281ff",
          2671 => x"0654b014",
          2672 => x"53727d70",
          2673 => x"81055f34",
          2674 => x"81177509",
          2675 => x"81057077",
          2676 => x"079f2a51",
          2677 => x"5457769f",
          2678 => x"26853872",
          2679 => x"ffaf3879",
          2680 => x"842a7081",
          2681 => x"06515372",
          2682 => x"802e8e38",
          2683 => x"963d7705",
          2684 => x"e00553ad",
          2685 => x"73348117",
          2686 => x"57767a81",
          2687 => x"065455b0",
          2688 => x"54728338",
          2689 => x"a0547981",
          2690 => x"2a708106",
          2691 => x"5456729f",
          2692 => x"38811755",
          2693 => x"767b2797",
          2694 => x"387351f9",
          2695 => x"f13f7581",
          2696 => x"0653728b",
          2697 => x"38748116",
          2698 => x"56537a73",
          2699 => x"26eb3896",
          2700 => x"3d7705e0",
          2701 => x"0553ff17",
          2702 => x"ff147033",
          2703 => x"535457f9",
          2704 => x"cd3f76f2",
          2705 => x"38748116",
          2706 => x"5653727b",
          2707 => x"27faf838",
          2708 => x"a051f9ba",
          2709 => x"3fef3996",
          2710 => x"3d0d04fd",
          2711 => x"3d0d863d",
          2712 => x"70708405",
          2713 => x"52085552",
          2714 => x"7351fad4",
          2715 => x"3f853d0d",
          2716 => x"04fe3d0d",
          2717 => x"74829cfc",
          2718 => x"0c853d88",
          2719 => x"05527551",
          2720 => x"fabe3f82",
          2721 => x"9cfc0853",
          2722 => x"80733480",
          2723 => x"0b829cfc",
          2724 => x"0c843d0d",
          2725 => x"04fd3d0d",
          2726 => x"829cf408",
          2727 => x"76829cf4",
          2728 => x"0c873d88",
          2729 => x"05537752",
          2730 => x"53fa953f",
          2731 => x"72829cf4",
          2732 => x"0c853d0d",
          2733 => x"04fb3d0d",
          2734 => x"7779829c",
          2735 => x"f8087056",
          2736 => x"54575580",
          2737 => x"5471802e",
          2738 => x"80e33882",
          2739 => x"9cf80852",
          2740 => x"712d8285",
          2741 => x"ec0881ff",
          2742 => x"06537280",
          2743 => x"2e80ce38",
          2744 => x"728d2ebc",
          2745 => x"38728832",
          2746 => x"70098105",
          2747 => x"70802551",
          2748 => x"51527380",
          2749 => x"2e8b3871",
          2750 => x"802e8638",
          2751 => x"ff145498",
          2752 => x"399f7325",
          2753 => x"c638ff16",
          2754 => x"52737225",
          2755 => x"ffbd3874",
          2756 => x"14527272",
          2757 => x"34811454",
          2758 => x"7251f7f2",
          2759 => x"3fffac39",
          2760 => x"73155280",
          2761 => x"72348a51",
          2762 => x"f7e43f81",
          2763 => x"53728285",
          2764 => x"ec0c873d",
          2765 => x"0d04fe3d",
          2766 => x"0d829cf8",
          2767 => x"0875829c",
          2768 => x"f80c7753",
          2769 => x"765253fe",
          2770 => x"ec3f7282",
          2771 => x"9cf80c84",
          2772 => x"3d0d04f8",
          2773 => x"3d0d7a7c",
          2774 => x"5a568070",
          2775 => x"7a0c5875",
          2776 => x"08703355",
          2777 => x"5373a02e",
          2778 => x"09810687",
          2779 => x"38811376",
          2780 => x"0ced3973",
          2781 => x"ad2e0981",
          2782 => x"068e3881",
          2783 => x"76081177",
          2784 => x"0c760870",
          2785 => x"33565458",
          2786 => x"73b02e09",
          2787 => x"810680c2",
          2788 => x"38750881",
          2789 => x"05760c75",
          2790 => x"08703355",
          2791 => x"537380e2",
          2792 => x"2e8b3890",
          2793 => x"577380f8",
          2794 => x"2e85388f",
          2795 => x"39825781",
          2796 => x"13760c75",
          2797 => x"08703355",
          2798 => x"53ac3981",
          2799 => x"55a07427",
          2800 => x"818438d0",
          2801 => x"14538055",
          2802 => x"88578973",
          2803 => x"27983880",
          2804 => x"f539d014",
          2805 => x"53805572",
          2806 => x"892680ea",
          2807 => x"38863980",
          2808 => x"5580e339",
          2809 => x"8a578055",
          2810 => x"a0742780",
          2811 => x"ca3880e0",
          2812 => x"74278938",
          2813 => x"e0147081",
          2814 => x"ff065553",
          2815 => x"d0147081",
          2816 => x"ff065553",
          2817 => x"9074278e",
          2818 => x"38f91470",
          2819 => x"81ff0655",
          2820 => x"53897427",
          2821 => x"ca387377",
          2822 => x"27c53876",
          2823 => x"527451c4",
          2824 => x"e93f8285",
          2825 => x"ec081476",
          2826 => x"08810577",
          2827 => x"0c760870",
          2828 => x"33565455",
          2829 => x"ffb23977",
          2830 => x"802e8638",
          2831 => x"74098105",
          2832 => x"5574790c",
          2833 => x"81557482",
          2834 => x"85ec0c8a",
          2835 => x"3d0d04f8",
          2836 => x"3d0d7a7c",
          2837 => x"5a568070",
          2838 => x"7a0c5875",
          2839 => x"08703355",
          2840 => x"5373a02e",
          2841 => x"09810687",
          2842 => x"38811376",
          2843 => x"0ced3973",
          2844 => x"ad2e0981",
          2845 => x"068e3881",
          2846 => x"76081177",
          2847 => x"0c760870",
          2848 => x"33565458",
          2849 => x"73b02e09",
          2850 => x"810680c2",
          2851 => x"38750881",
          2852 => x"05760c75",
          2853 => x"08703355",
          2854 => x"537380e2",
          2855 => x"2e8b3890",
          2856 => x"577380f8",
          2857 => x"2e85388f",
          2858 => x"39825781",
          2859 => x"13760c75",
          2860 => x"08703355",
          2861 => x"53ac3981",
          2862 => x"55a07427",
          2863 => x"818438d0",
          2864 => x"14538055",
          2865 => x"88578973",
          2866 => x"27983880",
          2867 => x"f539d014",
          2868 => x"53805572",
          2869 => x"892680ea",
          2870 => x"38863980",
          2871 => x"5580e339",
          2872 => x"8a578055",
          2873 => x"a0742780",
          2874 => x"ca3880e0",
          2875 => x"74278938",
          2876 => x"e0147081",
          2877 => x"ff065553",
          2878 => x"d0147081",
          2879 => x"ff065553",
          2880 => x"9074278e",
          2881 => x"38f91470",
          2882 => x"81ff0655",
          2883 => x"53897427",
          2884 => x"ca387377",
          2885 => x"27c53876",
          2886 => x"527451c2",
          2887 => x"ed3f8285",
          2888 => x"ec081476",
          2889 => x"08810577",
          2890 => x"0c760870",
          2891 => x"33565455",
          2892 => x"ffb23977",
          2893 => x"802e8638",
          2894 => x"74098105",
          2895 => x"5574790c",
          2896 => x"81557482",
          2897 => x"85ec0c8a",
          2898 => x"3d0d04fd",
          2899 => x"3d0d7698",
          2900 => x"2b70982c",
          2901 => x"79982b70",
          2902 => x"982c7210",
          2903 => x"7311822b",
          2904 => x"54565155",
          2905 => x"5151800b",
          2906 => x"81faf812",
          2907 => x"33555272",
          2908 => x"7425a038",
          2909 => x"7181faf4",
          2910 => x"12081402",
          2911 => x"88059705",
          2912 => x"33713352",
          2913 => x"53535470",
          2914 => x"722e0981",
          2915 => x"06833881",
          2916 => x"54735271",
          2917 => x"8285ec0c",
          2918 => x"853d0d04",
          2919 => x"fc3d0d78",
          2920 => x"0284059f",
          2921 => x"05337133",
          2922 => x"54555371",
          2923 => x"802e9f38",
          2924 => x"8851f2da",
          2925 => x"3fa051f2",
          2926 => x"d53f8851",
          2927 => x"f2d03f72",
          2928 => x"33ff0552",
          2929 => x"71733471",
          2930 => x"81ff0652",
          2931 => x"de397651",
          2932 => x"f3993f73",
          2933 => x"7334863d",
          2934 => x"0d04f63d",
          2935 => x"0d7c0284",
          2936 => x"05b70533",
          2937 => x"028805bb",
          2938 => x"05338285",
          2939 => x"c4337082",
          2940 => x"2b8284ec",
          2941 => x"11085159",
          2942 => x"595a5859",
          2943 => x"74802e86",
          2944 => x"3874519a",
          2945 => x"873f8285",
          2946 => x"c4337082",
          2947 => x"2b8284ec",
          2948 => x"11811a70",
          2949 => x"55595156",
          2950 => x"5a9d883f",
          2951 => x"8285ec08",
          2952 => x"750c8285",
          2953 => x"c4337082",
          2954 => x"2b8284ec",
          2955 => x"11085156",
          2956 => x"5a74802e",
          2957 => x"a7387553",
          2958 => x"78527451",
          2959 => x"ffb8da3f",
          2960 => x"8285c433",
          2961 => x"81055574",
          2962 => x"8285c434",
          2963 => x"7481ff06",
          2964 => x"55937527",
          2965 => x"8738800b",
          2966 => x"8285c434",
          2967 => x"77802eb6",
          2968 => x"388285c0",
          2969 => x"08567580",
          2970 => x"2eac3882",
          2971 => x"85bc3355",
          2972 => x"74a4388c",
          2973 => x"3dfc0554",
          2974 => x"76537852",
          2975 => x"755180d5",
          2976 => x"9f3f8285",
          2977 => x"c008528a",
          2978 => x"51818acd",
          2979 => x"3f8285c0",
          2980 => x"085180d8",
          2981 => x"fc3f8c3d",
          2982 => x"0d04fd3d",
          2983 => x"0d8284ec",
          2984 => x"53935472",
          2985 => x"08527180",
          2986 => x"2e893871",
          2987 => x"5198dd3f",
          2988 => x"80730cff",
          2989 => x"14841454",
          2990 => x"54738025",
          2991 => x"e638800b",
          2992 => x"8285c434",
          2993 => x"8285c008",
          2994 => x"5271802e",
          2995 => x"95387151",
          2996 => x"80d9dc3f",
          2997 => x"8285c008",
          2998 => x"5198b13f",
          2999 => x"800b8285",
          3000 => x"c00c853d",
          3001 => x"0d04dc3d",
          3002 => x"0d815780",
          3003 => x"528285c0",
          3004 => x"085180de",
          3005 => x"c83f8285",
          3006 => x"ec0880d2",
          3007 => x"388285c0",
          3008 => x"085380f8",
          3009 => x"52883d70",
          3010 => x"52568187",
          3011 => x"b33f8285",
          3012 => x"ec08802e",
          3013 => x"b9387551",
          3014 => x"ffb59e3f",
          3015 => x"8285ec08",
          3016 => x"55800b82",
          3017 => x"85ec0825",
          3018 => x"9c388285",
          3019 => x"ec08ff05",
          3020 => x"70175555",
          3021 => x"80743475",
          3022 => x"53765281",
          3023 => x"1781fde8",
          3024 => x"5257f697",
          3025 => x"3f74ff2e",
          3026 => x"098106ff",
          3027 => x"b038a63d",
          3028 => x"0d04d93d",
          3029 => x"0daa3d08",
          3030 => x"ad3d085a",
          3031 => x"5a817058",
          3032 => x"58805282",
          3033 => x"85c00851",
          3034 => x"80ddd23f",
          3035 => x"8285ec08",
          3036 => x"819638ff",
          3037 => x"0b8285c0",
          3038 => x"08545580",
          3039 => x"f8528b3d",
          3040 => x"70525681",
          3041 => x"86ba3f82",
          3042 => x"85ec0880",
          3043 => x"2ea53875",
          3044 => x"51ffb4a5",
          3045 => x"3f8285ec",
          3046 => x"08811858",
          3047 => x"55800b82",
          3048 => x"85ec0825",
          3049 => x"8e388285",
          3050 => x"ec08ff05",
          3051 => x"70175555",
          3052 => x"80743474",
          3053 => x"09700981",
          3054 => x"05707207",
          3055 => x"9f2a5155",
          3056 => x"5578772e",
          3057 => x"853873ff",
          3058 => x"aa388285",
          3059 => x"c0088c11",
          3060 => x"08535180",
          3061 => x"dce73f82",
          3062 => x"85ec0880",
          3063 => x"2e883881",
          3064 => x"fdf451ef",
          3065 => x"863f7877",
          3066 => x"2e098106",
          3067 => x"9b387552",
          3068 => x"7951ffb4",
          3069 => x"b23f7951",
          3070 => x"ffb3be3f",
          3071 => x"ab3d0854",
          3072 => x"8285ec08",
          3073 => x"74348058",
          3074 => x"778285ec",
          3075 => x"0ca93d0d",
          3076 => x"04f63d0d",
          3077 => x"7c7e715c",
          3078 => x"71723357",
          3079 => x"595a5873",
          3080 => x"a02e0981",
          3081 => x"06a23878",
          3082 => x"33780556",
          3083 => x"77762798",
          3084 => x"38811770",
          3085 => x"5b707133",
          3086 => x"56585573",
          3087 => x"a02e0981",
          3088 => x"06863875",
          3089 => x"7526ea38",
          3090 => x"80557483",
          3091 => x"2b8285c8",
          3092 => x"11700853",
          3093 => x"5154ffb2",
          3094 => x"e03f8285",
          3095 => x"ec085379",
          3096 => x"52730851",
          3097 => x"ffb5df3f",
          3098 => x"8285ec08",
          3099 => x"80c33884",
          3100 => x"14335473",
          3101 => x"812e8838",
          3102 => x"73822e88",
          3103 => x"38b339fc",
          3104 => x"e53fbe39",
          3105 => x"811a5a8c",
          3106 => x"3dfc1153",
          3107 => x"f80551f5",
          3108 => x"c23f8285",
          3109 => x"ec08802e",
          3110 => x"9838ff1b",
          3111 => x"53785277",
          3112 => x"51fdaf3f",
          3113 => x"8285ec08",
          3114 => x"81ff0654",
          3115 => x"73802e91",
          3116 => x"38811570",
          3117 => x"81ff0656",
          3118 => x"54827527",
          3119 => x"ff8c3880",
          3120 => x"54738285",
          3121 => x"ec0c8c3d",
          3122 => x"0d04d33d",
          3123 => x"0db03d08",
          3124 => x"b23d08b4",
          3125 => x"3d08595f",
          3126 => x"5a800baf",
          3127 => x"3d348285",
          3128 => x"c4338285",
          3129 => x"c008555b",
          3130 => x"7381ca38",
          3131 => x"738285bc",
          3132 => x"33555573",
          3133 => x"83388155",
          3134 => x"76802e81",
          3135 => x"bb388170",
          3136 => x"76065556",
          3137 => x"73802e81",
          3138 => x"ac38a851",
          3139 => x"97953f82",
          3140 => x"85ec0882",
          3141 => x"85c00c82",
          3142 => x"85ec0880",
          3143 => x"2e819138",
          3144 => x"93537652",
          3145 => x"8285ec08",
          3146 => x"5180c890",
          3147 => x"3f8285ec",
          3148 => x"08802e8b",
          3149 => x"3881fea0",
          3150 => x"51f2a03f",
          3151 => x"80f73982",
          3152 => x"85ec085b",
          3153 => x"8285c008",
          3154 => x"5380f852",
          3155 => x"903d7052",
          3156 => x"548182ec",
          3157 => x"3f8285ec",
          3158 => x"08568285",
          3159 => x"ec08742e",
          3160 => x"09810680",
          3161 => x"d0388285",
          3162 => x"ec0851ff",
          3163 => x"b0cb3f82",
          3164 => x"85ec0855",
          3165 => x"800b8285",
          3166 => x"ec0825a9",
          3167 => x"388285ec",
          3168 => x"08ff0570",
          3169 => x"17555580",
          3170 => x"74348053",
          3171 => x"7481ff06",
          3172 => x"527551f8",
          3173 => x"c53f811b",
          3174 => x"7081ff06",
          3175 => x"5c54937b",
          3176 => x"27833880",
          3177 => x"5b74ff2e",
          3178 => x"098106ff",
          3179 => x"97388639",
          3180 => x"758285bc",
          3181 => x"34768c38",
          3182 => x"8285c008",
          3183 => x"802e8438",
          3184 => x"f9d83f8f",
          3185 => x"3d5de09c",
          3186 => x"3f8285ec",
          3187 => x"08982b70",
          3188 => x"982c5159",
          3189 => x"78ff2eee",
          3190 => x"387881ff",
          3191 => x"06829d84",
          3192 => x"3370982b",
          3193 => x"70982c82",
          3194 => x"9d803370",
          3195 => x"982b7097",
          3196 => x"2c71982c",
          3197 => x"0570822b",
          3198 => x"81faf411",
          3199 => x"08157033",
          3200 => x"51515151",
          3201 => x"59595159",
          3202 => x"5d588156",
          3203 => x"73782e80",
          3204 => x"e3387774",
          3205 => x"27b138ff",
          3206 => x"1570982b",
          3207 => x"70982c51",
          3208 => x"56548075",
          3209 => x"2480cb38",
          3210 => x"76537452",
          3211 => x"7751f69b",
          3212 => x"3f8285ec",
          3213 => x"0881ff06",
          3214 => x"5473802e",
          3215 => x"da387482",
          3216 => x"9d803481",
          3217 => x"56ae3981",
          3218 => x"1570982b",
          3219 => x"70982c70",
          3220 => x"81ff0653",
          3221 => x"51565473",
          3222 => x"95269738",
          3223 => x"76537452",
          3224 => x"7751f5e7",
          3225 => x"3f8285ec",
          3226 => x"0881ff06",
          3227 => x"5473cf38",
          3228 => x"d6398056",
          3229 => x"75802e80",
          3230 => x"ca38811c",
          3231 => x"5473829d",
          3232 => x"84347398",
          3233 => x"2b70982c",
          3234 => x"829d8033",
          3235 => x"70982b70",
          3236 => x"982c7010",
          3237 => x"7111822b",
          3238 => x"81faf811",
          3239 => x"335e5253",
          3240 => x"51585851",
          3241 => x"5473772e",
          3242 => x"098106fe",
          3243 => x"993881fa",
          3244 => x"fc15087d",
          3245 => x"0c800b82",
          3246 => x"9d843480",
          3247 => x"0b829d80",
          3248 => x"34923975",
          3249 => x"829d8434",
          3250 => x"75829d80",
          3251 => x"3478af3d",
          3252 => x"34757d0c",
          3253 => x"7e547395",
          3254 => x"26fde838",
          3255 => x"73822b54",
          3256 => x"81e8f014",
          3257 => x"0804829d",
          3258 => x"8c335675",
          3259 => x"7e2efdd3",
          3260 => x"38829d88",
          3261 => x"33547574",
          3262 => x"27ab3873",
          3263 => x"982b7098",
          3264 => x"2c515575",
          3265 => x"75249e38",
          3266 => x"741a5473",
          3267 => x"33811534",
          3268 => x"ff157098",
          3269 => x"2b70982c",
          3270 => x"829d8c33",
          3271 => x"53515654",
          3272 => x"747425e4",
          3273 => x"38829d8c",
          3274 => x"33811156",
          3275 => x"5474829d",
          3276 => x"8c34731a",
          3277 => x"54ae3d33",
          3278 => x"7434829d",
          3279 => x"88335473",
          3280 => x"7e258938",
          3281 => x"81145473",
          3282 => x"829d8834",
          3283 => x"829d8c33",
          3284 => x"ff057098",
          3285 => x"2b70982c",
          3286 => x"829d8833",
          3287 => x"59515654",
          3288 => x"7476259f",
          3289 => x"38741a70",
          3290 => x"335254e7",
          3291 => x"a13f8115",
          3292 => x"70982b70",
          3293 => x"982c829d",
          3294 => x"88335a51",
          3295 => x"56547675",
          3296 => x"24e33882",
          3297 => x"9d8c3370",
          3298 => x"982b7098",
          3299 => x"2c829d88",
          3300 => x"33595156",
          3301 => x"54747625",
          3302 => x"fca93888",
          3303 => x"51e6ef3f",
          3304 => x"81157098",
          3305 => x"2b70982c",
          3306 => x"829d8833",
          3307 => x"5a515654",
          3308 => x"767524e7",
          3309 => x"38fc8c39",
          3310 => x"837a3480",
          3311 => x"0b811b34",
          3312 => x"829d8c53",
          3313 => x"805281f3",
          3314 => x"d851f3d0",
          3315 => x"3f81d939",
          3316 => x"829d8c33",
          3317 => x"7081ff06",
          3318 => x"55557380",
          3319 => x"2efbe438",
          3320 => x"829d8833",
          3321 => x"ff055473",
          3322 => x"829d8834",
          3323 => x"ff155473",
          3324 => x"829d8c34",
          3325 => x"8851e696",
          3326 => x"3f829d8c",
          3327 => x"3370982b",
          3328 => x"70982c82",
          3329 => x"9d883357",
          3330 => x"51565774",
          3331 => x"7425a438",
          3332 => x"741a5481",
          3333 => x"14337434",
          3334 => x"733351e5",
          3335 => x"f13f8115",
          3336 => x"70982b70",
          3337 => x"982c829d",
          3338 => x"88335951",
          3339 => x"56547575",
          3340 => x"24de38a0",
          3341 => x"51e5d73f",
          3342 => x"829d8c33",
          3343 => x"70982b70",
          3344 => x"982c829d",
          3345 => x"88335751",
          3346 => x"56577474",
          3347 => x"24faf438",
          3348 => x"8851e5ba",
          3349 => x"3f811570",
          3350 => x"982b7098",
          3351 => x"2c829d88",
          3352 => x"33595156",
          3353 => x"54757525",
          3354 => x"e738fad7",
          3355 => x"39829d88",
          3356 => x"337a0554",
          3357 => x"8074348a",
          3358 => x"51e5933f",
          3359 => x"829d8852",
          3360 => x"7951f78d",
          3361 => x"3f8285ec",
          3362 => x"0881ff06",
          3363 => x"54739638",
          3364 => x"829d8833",
          3365 => x"5473802e",
          3366 => x"8f388153",
          3367 => x"73527951",
          3368 => x"f2b83f84",
          3369 => x"39807a34",
          3370 => x"800b829d",
          3371 => x"8c34800b",
          3372 => x"829d8834",
          3373 => x"798285ec",
          3374 => x"0caf3d0d",
          3375 => x"04829d8c",
          3376 => x"33547380",
          3377 => x"2ef9fc38",
          3378 => x"8851e4c2",
          3379 => x"3f829d8c",
          3380 => x"33ff0554",
          3381 => x"73829d8c",
          3382 => x"347381ff",
          3383 => x"0654e339",
          3384 => x"829d8c33",
          3385 => x"829d8833",
          3386 => x"55557375",
          3387 => x"2ef9d438",
          3388 => x"ff145473",
          3389 => x"829d8834",
          3390 => x"74982b70",
          3391 => x"982c7581",
          3392 => x"ff065651",
          3393 => x"55747425",
          3394 => x"a438741a",
          3395 => x"54811433",
          3396 => x"74347333",
          3397 => x"51e3f73f",
          3398 => x"81157098",
          3399 => x"2b70982c",
          3400 => x"829d8833",
          3401 => x"59515654",
          3402 => x"757524de",
          3403 => x"38a051e3",
          3404 => x"dd3f829d",
          3405 => x"8c337098",
          3406 => x"2b70982c",
          3407 => x"829d8833",
          3408 => x"57515657",
          3409 => x"747424f8",
          3410 => x"fa388851",
          3411 => x"e3c03f81",
          3412 => x"1570982b",
          3413 => x"70982c82",
          3414 => x"9d883359",
          3415 => x"51565475",
          3416 => x"7525e738",
          3417 => x"f8dd3982",
          3418 => x"9d8c3370",
          3419 => x"81ff0682",
          3420 => x"9d883359",
          3421 => x"56547477",
          3422 => x"27f8c838",
          3423 => x"81145473",
          3424 => x"829d8c34",
          3425 => x"741a7033",
          3426 => x"5254e382",
          3427 => x"3f829d8c",
          3428 => x"337081ff",
          3429 => x"06829d88",
          3430 => x"33585654",
          3431 => x"757526dc",
          3432 => x"38f8a039",
          3433 => x"829d8c53",
          3434 => x"805281f3",
          3435 => x"d851efec",
          3436 => x"3f800b82",
          3437 => x"9d8c3480",
          3438 => x"0b829d88",
          3439 => x"34f88439",
          3440 => x"7ab03882",
          3441 => x"85b80855",
          3442 => x"74802ea6",
          3443 => x"387451ff",
          3444 => x"a7e73f82",
          3445 => x"85ec0882",
          3446 => x"9d883482",
          3447 => x"85ec0881",
          3448 => x"ff068105",
          3449 => x"53745279",
          3450 => x"51ffa9ad",
          3451 => x"3f935b81",
          3452 => x"c0397a82",
          3453 => x"2b8284ec",
          3454 => x"11fc1108",
          3455 => x"57515474",
          3456 => x"802ea738",
          3457 => x"7451ffa7",
          3458 => x"b03f8285",
          3459 => x"ec08829d",
          3460 => x"88348285",
          3461 => x"ec0881ff",
          3462 => x"06810553",
          3463 => x"74527951",
          3464 => x"ffa8f63f",
          3465 => x"ff1b5480",
          3466 => x"f9397308",
          3467 => x"5574802e",
          3468 => x"f7913874",
          3469 => x"51ffa781",
          3470 => x"3f99397a",
          3471 => x"932e0981",
          3472 => x"06ae3882",
          3473 => x"84ec0855",
          3474 => x"74802ea4",
          3475 => x"387451ff",
          3476 => x"a6e73f82",
          3477 => x"85ec0882",
          3478 => x"9d883482",
          3479 => x"85ec0881",
          3480 => x"ff068105",
          3481 => x"53745279",
          3482 => x"51ffa8ad",
          3483 => x"3f80c239",
          3484 => x"7a822b82",
          3485 => x"84f01108",
          3486 => x"56547480",
          3487 => x"2eab3874",
          3488 => x"51ffa6b5",
          3489 => x"3f8285ec",
          3490 => x"08829d88",
          3491 => x"348285ec",
          3492 => x"0881ff06",
          3493 => x"81055374",
          3494 => x"527951ff",
          3495 => x"a7fb3f81",
          3496 => x"1b547381",
          3497 => x"ff065b89",
          3498 => x"3974829d",
          3499 => x"8834747a",
          3500 => x"34829d8c",
          3501 => x"53829d88",
          3502 => x"33527951",
          3503 => x"edde3ff6",
          3504 => x"8239829d",
          3505 => x"8c337081",
          3506 => x"ff06829d",
          3507 => x"88335956",
          3508 => x"54747727",
          3509 => x"f5ed3881",
          3510 => x"14547382",
          3511 => x"9d8c3474",
          3512 => x"1a703352",
          3513 => x"54e0a73f",
          3514 => x"f5d93982",
          3515 => x"9d8c3354",
          3516 => x"73802ef5",
          3517 => x"ce388851",
          3518 => x"e0943f82",
          3519 => x"9d8c33ff",
          3520 => x"05547382",
          3521 => x"9d8c34f5",
          3522 => x"ba39f93d",
          3523 => x"0d83dff4",
          3524 => x"0b8285e4",
          3525 => x"0c82800b",
          3526 => x"8285e023",
          3527 => x"90805380",
          3528 => x"5283dff4",
          3529 => x"51ffaac5",
          3530 => x"3f8285e4",
          3531 => x"08548058",
          3532 => x"77743481",
          3533 => x"57768115",
          3534 => x"348285e4",
          3535 => x"08547784",
          3536 => x"15347685",
          3537 => x"15348285",
          3538 => x"e4085477",
          3539 => x"86153476",
          3540 => x"87153482",
          3541 => x"85e40882",
          3542 => x"85e022ff",
          3543 => x"05fe8080",
          3544 => x"077083ff",
          3545 => x"ff067088",
          3546 => x"2a585155",
          3547 => x"56748817",
          3548 => x"34738917",
          3549 => x"348285e0",
          3550 => x"2270832b",
          3551 => x"8285e408",
          3552 => x"11f80551",
          3553 => x"55557782",
          3554 => x"15347683",
          3555 => x"1534893d",
          3556 => x"0d04ff3d",
          3557 => x"0d735281",
          3558 => x"51847227",
          3559 => x"8f38fb12",
          3560 => x"832a8211",
          3561 => x"7083ffff",
          3562 => x"06515151",
          3563 => x"708285ec",
          3564 => x"0c833d0d",
          3565 => x"04f93d0d",
          3566 => x"02a60522",
          3567 => x"028405aa",
          3568 => x"05227105",
          3569 => x"8285e408",
          3570 => x"71832b71",
          3571 => x"1174832b",
          3572 => x"73117033",
          3573 => x"81123371",
          3574 => x"882b0702",
          3575 => x"a405ae05",
          3576 => x"227181ff",
          3577 => x"ff060770",
          3578 => x"882a5351",
          3579 => x"5259545b",
          3580 => x"5b575354",
          3581 => x"55717734",
          3582 => x"70811834",
          3583 => x"8285e408",
          3584 => x"1475882a",
          3585 => x"52547082",
          3586 => x"15347483",
          3587 => x"15348285",
          3588 => x"e4087017",
          3589 => x"70338112",
          3590 => x"3371882b",
          3591 => x"0770832b",
          3592 => x"8ffff806",
          3593 => x"51525652",
          3594 => x"71057383",
          3595 => x"ffff0670",
          3596 => x"882a5454",
          3597 => x"51718212",
          3598 => x"347281ff",
          3599 => x"06537283",
          3600 => x"12348285",
          3601 => x"e4081656",
          3602 => x"71763472",
          3603 => x"81173489",
          3604 => x"3d0d04fb",
          3605 => x"3d0d8285",
          3606 => x"e4080284",
          3607 => x"059e0522",
          3608 => x"70832b72",
          3609 => x"11861133",
          3610 => x"87123371",
          3611 => x"8b2b7183",
          3612 => x"2b07585b",
          3613 => x"59525552",
          3614 => x"72058412",
          3615 => x"33851333",
          3616 => x"71882b07",
          3617 => x"70882a54",
          3618 => x"56565270",
          3619 => x"84133473",
          3620 => x"85133482",
          3621 => x"85e40870",
          3622 => x"14841133",
          3623 => x"85123371",
          3624 => x"8b2b7183",
          3625 => x"2b075659",
          3626 => x"57527205",
          3627 => x"86123387",
          3628 => x"13337188",
          3629 => x"2b077088",
          3630 => x"2a545656",
          3631 => x"52708613",
          3632 => x"34738713",
          3633 => x"348285e4",
          3634 => x"08137033",
          3635 => x"81123371",
          3636 => x"882b0770",
          3637 => x"81ffff06",
          3638 => x"70882a53",
          3639 => x"51535353",
          3640 => x"71733470",
          3641 => x"81143487",
          3642 => x"3d0d04f9",
          3643 => x"3d0d02a6",
          3644 => x"05228285",
          3645 => x"e4087183",
          3646 => x"2b711170",
          3647 => x"33811233",
          3648 => x"71882b07",
          3649 => x"70832b53",
          3650 => x"595b5558",
          3651 => x"73057033",
          3652 => x"81123371",
          3653 => x"982b7190",
          3654 => x"2b07535a",
          3655 => x"55535571",
          3656 => x"802580f6",
          3657 => x"387351fe",
          3658 => x"aa3f8285",
          3659 => x"e4087017",
          3660 => x"70338112",
          3661 => x"33718b2b",
          3662 => x"71832b07",
          3663 => x"74117033",
          3664 => x"81123371",
          3665 => x"882b0770",
          3666 => x"832b8fff",
          3667 => x"f8065152",
          3668 => x"5d515357",
          3669 => x"5a537205",
          3670 => x"75882a54",
          3671 => x"52728213",
          3672 => x"34748313",
          3673 => x"348285e4",
          3674 => x"08701770",
          3675 => x"33811233",
          3676 => x"718b2b71",
          3677 => x"832b0756",
          3678 => x"59575572",
          3679 => x"05703381",
          3680 => x"12337188",
          3681 => x"2b077081",
          3682 => x"ffff0670",
          3683 => x"882a5751",
          3684 => x"52585272",
          3685 => x"74347181",
          3686 => x"1534893d",
          3687 => x"0d04fb3d",
          3688 => x"0d8285e4",
          3689 => x"08028405",
          3690 => x"9e052270",
          3691 => x"832b7211",
          3692 => x"82113383",
          3693 => x"1233718b",
          3694 => x"2b71832b",
          3695 => x"07595b59",
          3696 => x"52565273",
          3697 => x"05713381",
          3698 => x"13337188",
          3699 => x"2b07028c",
          3700 => x"05a20522",
          3701 => x"71077088",
          3702 => x"2a535153",
          3703 => x"53537173",
          3704 => x"34708114",
          3705 => x"348285e4",
          3706 => x"08701570",
          3707 => x"33811233",
          3708 => x"718b2b71",
          3709 => x"832b0756",
          3710 => x"59575272",
          3711 => x"05821233",
          3712 => x"83133371",
          3713 => x"882b0770",
          3714 => x"882a5455",
          3715 => x"56527082",
          3716 => x"13347283",
          3717 => x"13348285",
          3718 => x"e4081482",
          3719 => x"11338312",
          3720 => x"3371882b",
          3721 => x"078285ec",
          3722 => x"0c525487",
          3723 => x"3d0d04f7",
          3724 => x"3d0d7b82",
          3725 => x"85e40831",
          3726 => x"832a7083",
          3727 => x"ffff0670",
          3728 => x"535753fd",
          3729 => x"a63f8285",
          3730 => x"e4087683",
          3731 => x"2b711182",
          3732 => x"11338312",
          3733 => x"33718b2b",
          3734 => x"71832b07",
          3735 => x"75117033",
          3736 => x"81123371",
          3737 => x"982b7190",
          3738 => x"2b075342",
          3739 => x"4051535b",
          3740 => x"58555954",
          3741 => x"7280258d",
          3742 => x"38828080",
          3743 => x"527551fe",
          3744 => x"9d3f8184",
          3745 => x"39841433",
          3746 => x"85153371",
          3747 => x"8b2b7183",
          3748 => x"2b077611",
          3749 => x"79882a53",
          3750 => x"51555855",
          3751 => x"76861434",
          3752 => x"7581ff06",
          3753 => x"56758714",
          3754 => x"348285e4",
          3755 => x"08701984",
          3756 => x"12338513",
          3757 => x"3371882b",
          3758 => x"0770882a",
          3759 => x"54575b56",
          3760 => x"53728416",
          3761 => x"34738516",
          3762 => x"348285e4",
          3763 => x"08185380",
          3764 => x"0b861434",
          3765 => x"800b8714",
          3766 => x"348285e4",
          3767 => x"08537684",
          3768 => x"14347585",
          3769 => x"14348285",
          3770 => x"e4081870",
          3771 => x"33811233",
          3772 => x"71882b07",
          3773 => x"70828080",
          3774 => x"0770882a",
          3775 => x"53515556",
          3776 => x"54747434",
          3777 => x"72811534",
          3778 => x"8b3d0d04",
          3779 => x"ff3d0d73",
          3780 => x"528285e4",
          3781 => x"088438f7",
          3782 => x"f13f7180",
          3783 => x"2e863871",
          3784 => x"51fe8c3f",
          3785 => x"833d0d04",
          3786 => x"f53d0d80",
          3787 => x"7e5258f8",
          3788 => x"e13f8285",
          3789 => x"ec0883ff",
          3790 => x"ff068285",
          3791 => x"e4088411",
          3792 => x"33851233",
          3793 => x"71882b07",
          3794 => x"705f5956",
          3795 => x"585a81ff",
          3796 => x"ff597578",
          3797 => x"2e80cc38",
          3798 => x"75832b77",
          3799 => x"05703381",
          3800 => x"12337188",
          3801 => x"2b077081",
          3802 => x"ffff0679",
          3803 => x"317083ff",
          3804 => x"ff06707f",
          3805 => x"27525351",
          3806 => x"56595577",
          3807 => x"79278a38",
          3808 => x"73802e85",
          3809 => x"3875785a",
          3810 => x"5b841533",
          3811 => x"85163371",
          3812 => x"882b0757",
          3813 => x"5475c138",
          3814 => x"7881ffff",
          3815 => x"2e85387a",
          3816 => x"79595680",
          3817 => x"76832b82",
          3818 => x"85e40811",
          3819 => x"70338112",
          3820 => x"3371882b",
          3821 => x"077081ff",
          3822 => x"ff065152",
          3823 => x"5a565c55",
          3824 => x"73752e83",
          3825 => x"38815580",
          3826 => x"54797826",
          3827 => x"81cc3874",
          3828 => x"5474802e",
          3829 => x"81c43877",
          3830 => x"7a2e0981",
          3831 => x"06893875",
          3832 => x"51f8f03f",
          3833 => x"81ac3982",
          3834 => x"80805379",
          3835 => x"527551f7",
          3836 => x"c43f8285",
          3837 => x"e408701c",
          3838 => x"86113387",
          3839 => x"1233718b",
          3840 => x"2b71832b",
          3841 => x"07535a5e",
          3842 => x"5574057a",
          3843 => x"177083ff",
          3844 => x"ff067088",
          3845 => x"2a5c5956",
          3846 => x"54788415",
          3847 => x"347681ff",
          3848 => x"06577685",
          3849 => x"15348285",
          3850 => x"e4087583",
          3851 => x"2b711172",
          3852 => x"1e861133",
          3853 => x"87123371",
          3854 => x"882b0770",
          3855 => x"882a535b",
          3856 => x"5e535a56",
          3857 => x"54738619",
          3858 => x"34758719",
          3859 => x"348285e4",
          3860 => x"08701c84",
          3861 => x"11338512",
          3862 => x"33718b2b",
          3863 => x"71832b07",
          3864 => x"535d5a55",
          3865 => x"74055478",
          3866 => x"86153476",
          3867 => x"87153482",
          3868 => x"85e40870",
          3869 => x"16711d84",
          3870 => x"11338512",
          3871 => x"3371882b",
          3872 => x"0770882a",
          3873 => x"535a5f52",
          3874 => x"56547384",
          3875 => x"16347585",
          3876 => x"16348285",
          3877 => x"e4081b84",
          3878 => x"05547382",
          3879 => x"85ec0c8d",
          3880 => x"3d0d04fe",
          3881 => x"3d0d7452",
          3882 => x"8285e408",
          3883 => x"8438f4da",
          3884 => x"3f715371",
          3885 => x"802e8b38",
          3886 => x"7151fcec",
          3887 => x"3f8285ec",
          3888 => x"08537282",
          3889 => x"85ec0c84",
          3890 => x"3d0d04ff",
          3891 => x"3d0d028f",
          3892 => x"05335181",
          3893 => x"52707226",
          3894 => x"87388285",
          3895 => x"e8113352",
          3896 => x"718285ec",
          3897 => x"0c833d0d",
          3898 => x"04fc3d0d",
          3899 => x"029b0533",
          3900 => x"0284059f",
          3901 => x"05335653",
          3902 => x"83517281",
          3903 => x"2680e038",
          3904 => x"72842b87",
          3905 => x"c0928c11",
          3906 => x"53518854",
          3907 => x"74802e84",
          3908 => x"38818854",
          3909 => x"73720c87",
          3910 => x"c0928c11",
          3911 => x"5181710c",
          3912 => x"850b87c0",
          3913 => x"988c0c70",
          3914 => x"52710870",
          3915 => x"82065151",
          3916 => x"70802e8a",
          3917 => x"3887c098",
          3918 => x"8c085170",
          3919 => x"ec387108",
          3920 => x"fc808006",
          3921 => x"52719238",
          3922 => x"87c0988c",
          3923 => x"08517080",
          3924 => x"2e873871",
          3925 => x"8285e814",
          3926 => x"348285e8",
          3927 => x"13335170",
          3928 => x"8285ec0c",
          3929 => x"863d0d04",
          3930 => x"f33d0d60",
          3931 => x"6264028c",
          3932 => x"05bf0533",
          3933 => x"5740585b",
          3934 => x"8374525a",
          3935 => x"fecd3f82",
          3936 => x"85ec0881",
          3937 => x"067a5452",
          3938 => x"7181be38",
          3939 => x"71727584",
          3940 => x"2b87c092",
          3941 => x"801187c0",
          3942 => x"928c1287",
          3943 => x"c0928413",
          3944 => x"415a4057",
          3945 => x"5a58850b",
          3946 => x"87c0988c",
          3947 => x"0c767d0c",
          3948 => x"84760c75",
          3949 => x"0870852a",
          3950 => x"70810651",
          3951 => x"53547180",
          3952 => x"2e8e387b",
          3953 => x"0852717b",
          3954 => x"7081055d",
          3955 => x"34811959",
          3956 => x"8074a206",
          3957 => x"53537173",
          3958 => x"2e833881",
          3959 => x"537883ff",
          3960 => x"268f3872",
          3961 => x"802e8a38",
          3962 => x"87c0988c",
          3963 => x"085271c3",
          3964 => x"3887c098",
          3965 => x"8c085271",
          3966 => x"802e8738",
          3967 => x"7884802e",
          3968 => x"99388176",
          3969 => x"0c87c092",
          3970 => x"8c155372",
          3971 => x"08708206",
          3972 => x"515271f7",
          3973 => x"38ff1a5a",
          3974 => x"8d398480",
          3975 => x"17811970",
          3976 => x"81ff065a",
          3977 => x"53577980",
          3978 => x"2e903873",
          3979 => x"fc808006",
          3980 => x"52718738",
          3981 => x"7d7826fe",
          3982 => x"ed3873fc",
          3983 => x"80800652",
          3984 => x"71802e83",
          3985 => x"38815271",
          3986 => x"53728285",
          3987 => x"ec0c8f3d",
          3988 => x"0d04f33d",
          3989 => x"0d606264",
          3990 => x"028c05bf",
          3991 => x"05335740",
          3992 => x"585b8359",
          3993 => x"80745258",
          3994 => x"fce13f82",
          3995 => x"85ec0881",
          3996 => x"06795452",
          3997 => x"71782e09",
          3998 => x"810681b1",
          3999 => x"38777484",
          4000 => x"2b87c092",
          4001 => x"801187c0",
          4002 => x"928c1287",
          4003 => x"c0928413",
          4004 => x"40595f56",
          4005 => x"5a850b87",
          4006 => x"c0988c0c",
          4007 => x"767d0c82",
          4008 => x"760c8058",
          4009 => x"75087084",
          4010 => x"2a708106",
          4011 => x"51535471",
          4012 => x"802e8c38",
          4013 => x"7a708105",
          4014 => x"5c337c0c",
          4015 => x"81185873",
          4016 => x"812a7081",
          4017 => x"06515271",
          4018 => x"802e8a38",
          4019 => x"87c0988c",
          4020 => x"085271d0",
          4021 => x"3887c098",
          4022 => x"8c085271",
          4023 => x"802e8738",
          4024 => x"7784802e",
          4025 => x"99388176",
          4026 => x"0c87c092",
          4027 => x"8c155372",
          4028 => x"08708206",
          4029 => x"515271f7",
          4030 => x"38ff1959",
          4031 => x"8d39811a",
          4032 => x"7081ff06",
          4033 => x"84801959",
          4034 => x"5b527880",
          4035 => x"2e903873",
          4036 => x"fc808006",
          4037 => x"52718738",
          4038 => x"7d7a26fe",
          4039 => x"f83873fc",
          4040 => x"80800652",
          4041 => x"71802e83",
          4042 => x"38815271",
          4043 => x"53728285",
          4044 => x"ec0c8f3d",
          4045 => x"0d04fa3d",
          4046 => x"0d7a0284",
          4047 => x"05a30533",
          4048 => x"028805a7",
          4049 => x"05337154",
          4050 => x"545657fa",
          4051 => x"fe3f8285",
          4052 => x"ec088106",
          4053 => x"53835472",
          4054 => x"80fe3885",
          4055 => x"0b87c098",
          4056 => x"8c0c8156",
          4057 => x"71762e80",
          4058 => x"dc387176",
          4059 => x"24933874",
          4060 => x"842b87c0",
          4061 => x"928c1154",
          4062 => x"5471802e",
          4063 => x"8d3880d4",
          4064 => x"3971832e",
          4065 => x"80c63880",
          4066 => x"cb397208",
          4067 => x"70812a70",
          4068 => x"81065151",
          4069 => x"5271802e",
          4070 => x"8a3887c0",
          4071 => x"988c0852",
          4072 => x"71e83887",
          4073 => x"c0988c08",
          4074 => x"52719638",
          4075 => x"81730c87",
          4076 => x"c0928c14",
          4077 => x"53720870",
          4078 => x"82065152",
          4079 => x"71f73896",
          4080 => x"39805692",
          4081 => x"3988800a",
          4082 => x"770c8539",
          4083 => x"8180770c",
          4084 => x"72568339",
          4085 => x"84567554",
          4086 => x"738285ec",
          4087 => x"0c883d0d",
          4088 => x"04fe3d0d",
          4089 => x"74811133",
          4090 => x"71337188",
          4091 => x"2b078285",
          4092 => x"ec0c5351",
          4093 => x"843d0d04",
          4094 => x"fd3d0d75",
          4095 => x"83113382",
          4096 => x"12337190",
          4097 => x"2b71882b",
          4098 => x"07811433",
          4099 => x"70720788",
          4100 => x"2b753371",
          4101 => x"078285ec",
          4102 => x"0c525354",
          4103 => x"56545285",
          4104 => x"3d0d04ff",
          4105 => x"3d0d7302",
          4106 => x"84059205",
          4107 => x"22525270",
          4108 => x"72708105",
          4109 => x"54347088",
          4110 => x"2a517072",
          4111 => x"34833d0d",
          4112 => x"04ff3d0d",
          4113 => x"73755252",
          4114 => x"70727081",
          4115 => x"05543470",
          4116 => x"882a5170",
          4117 => x"72708105",
          4118 => x"54347088",
          4119 => x"2a517072",
          4120 => x"70810554",
          4121 => x"3470882a",
          4122 => x"51707234",
          4123 => x"833d0d04",
          4124 => x"fe3d0d76",
          4125 => x"75775454",
          4126 => x"5170802e",
          4127 => x"92387170",
          4128 => x"81055333",
          4129 => x"73708105",
          4130 => x"5534ff11",
          4131 => x"51eb3984",
          4132 => x"3d0d04fe",
          4133 => x"3d0d7577",
          4134 => x"76545253",
          4135 => x"72727081",
          4136 => x"055434ff",
          4137 => x"115170f4",
          4138 => x"38843d0d",
          4139 => x"04fc3d0d",
          4140 => x"78777956",
          4141 => x"56537470",
          4142 => x"81055633",
          4143 => x"74708105",
          4144 => x"56337171",
          4145 => x"31ff1656",
          4146 => x"52525272",
          4147 => x"802e8638",
          4148 => x"71802ee2",
          4149 => x"38718285",
          4150 => x"ec0c863d",
          4151 => x"0d04fe3d",
          4152 => x"0d747654",
          4153 => x"51893971",
          4154 => x"732e8a38",
          4155 => x"81115170",
          4156 => x"335271f3",
          4157 => x"38703382",
          4158 => x"85ec0c84",
          4159 => x"3d0d0480",
          4160 => x"0b8285ec",
          4161 => x"0c04800b",
          4162 => x"8285ec0c",
          4163 => x"04f73d0d",
          4164 => x"7b56800b",
          4165 => x"83173356",
          4166 => x"5a747a2e",
          4167 => x"80d63881",
          4168 => x"54b01608",
          4169 => x"53b41670",
          4170 => x"53811733",
          4171 => x"5259faa2",
          4172 => x"3f8285ec",
          4173 => x"087a2e09",
          4174 => x"8106b738",
          4175 => x"8285ec08",
          4176 => x"831734b0",
          4177 => x"160870a4",
          4178 => x"1808319c",
          4179 => x"18085956",
          4180 => x"58747727",
          4181 => x"9f388216",
          4182 => x"33557482",
          4183 => x"2e098106",
          4184 => x"93388154",
          4185 => x"76185378",
          4186 => x"52811633",
          4187 => x"51f9e33f",
          4188 => x"8339815a",
          4189 => x"798285ec",
          4190 => x"0c8b3d0d",
          4191 => x"04fa3d0d",
          4192 => x"787a5656",
          4193 => x"805774b0",
          4194 => x"17082eaf",
          4195 => x"387551fe",
          4196 => x"fc3f8285",
          4197 => x"ec085782",
          4198 => x"85ec089f",
          4199 => x"38815474",
          4200 => x"53b41652",
          4201 => x"81163351",
          4202 => x"f7be3f82",
          4203 => x"85ec0880",
          4204 => x"2e8538ff",
          4205 => x"55815774",
          4206 => x"b0170c76",
          4207 => x"8285ec0c",
          4208 => x"883d0d04",
          4209 => x"f83d0d7a",
          4210 => x"705257fe",
          4211 => x"c03f8285",
          4212 => x"ec085882",
          4213 => x"85ec0881",
          4214 => x"91387633",
          4215 => x"5574832e",
          4216 => x"09810680",
          4217 => x"f0388417",
          4218 => x"33597881",
          4219 => x"2e098106",
          4220 => x"80e33884",
          4221 => x"80538285",
          4222 => x"ec0852b4",
          4223 => x"17705256",
          4224 => x"fd913f82",
          4225 => x"d4d55284",
          4226 => x"b21751fc",
          4227 => x"963f848b",
          4228 => x"85a4d252",
          4229 => x"7551fca9",
          4230 => x"3f868a85",
          4231 => x"e4f25284",
          4232 => x"981751fc",
          4233 => x"9c3f9017",
          4234 => x"0852849c",
          4235 => x"1751fc91",
          4236 => x"3f8c1708",
          4237 => x"5284a017",
          4238 => x"51fc863f",
          4239 => x"a0170881",
          4240 => x"0570b019",
          4241 => x"0c795553",
          4242 => x"75528117",
          4243 => x"3351f882",
          4244 => x"3f778418",
          4245 => x"34805380",
          4246 => x"52811733",
          4247 => x"51f9d73f",
          4248 => x"8285ec08",
          4249 => x"802e8338",
          4250 => x"81587782",
          4251 => x"85ec0c8a",
          4252 => x"3d0d04fb",
          4253 => x"3d0d77fe",
          4254 => x"1a981208",
          4255 => x"fe055555",
          4256 => x"55805673",
          4257 => x"73279438",
          4258 => x"8a152274",
          4259 => x"5351ff97",
          4260 => x"f93fac15",
          4261 => x"088285ec",
          4262 => x"08055675",
          4263 => x"8285ec0c",
          4264 => x"873d0d04",
          4265 => x"f93d0d7a",
          4266 => x"7a700856",
          4267 => x"54578177",
          4268 => x"2781df38",
          4269 => x"76981508",
          4270 => x"2781d738",
          4271 => x"ff743354",
          4272 => x"5872822e",
          4273 => x"80f53872",
          4274 => x"82248938",
          4275 => x"72812e8d",
          4276 => x"3881bf39",
          4277 => x"72832e81",
          4278 => x"8e3881b6",
          4279 => x"3976812a",
          4280 => x"1770892a",
          4281 => x"a4160805",
          4282 => x"53745255",
          4283 => x"fd8f3f82",
          4284 => x"85ec0881",
          4285 => x"9f387483",
          4286 => x"ff0614b4",
          4287 => x"11338117",
          4288 => x"70892aa4",
          4289 => x"18080555",
          4290 => x"76545757",
          4291 => x"53fcee3f",
          4292 => x"8285ec08",
          4293 => x"80fe3874",
          4294 => x"83ff0614",
          4295 => x"b4113370",
          4296 => x"882b7807",
          4297 => x"79810671",
          4298 => x"842a5c52",
          4299 => x"58515372",
          4300 => x"80e23875",
          4301 => x"9fff0658",
          4302 => x"80da3976",
          4303 => x"882aa415",
          4304 => x"08055273",
          4305 => x"51fcb63f",
          4306 => x"8285ec08",
          4307 => x"80c63876",
          4308 => x"1083fe06",
          4309 => x"7405b405",
          4310 => x"51f9863f",
          4311 => x"8285ec08",
          4312 => x"83ffff06",
          4313 => x"58ae3976",
          4314 => x"872aa415",
          4315 => x"08055273",
          4316 => x"51fc8a3f",
          4317 => x"8285ec08",
          4318 => x"9b387682",
          4319 => x"2b83fc06",
          4320 => x"7405b405",
          4321 => x"51f8f13f",
          4322 => x"8285ec08",
          4323 => x"f00a0658",
          4324 => x"83398158",
          4325 => x"778285ec",
          4326 => x"0c893d0d",
          4327 => x"04f83d0d",
          4328 => x"7a7c7e5a",
          4329 => x"58568259",
          4330 => x"81772782",
          4331 => x"9e387698",
          4332 => x"17082782",
          4333 => x"96387533",
          4334 => x"5372792e",
          4335 => x"819d3872",
          4336 => x"79248938",
          4337 => x"72812e8d",
          4338 => x"38828039",
          4339 => x"72832e81",
          4340 => x"b83881f7",
          4341 => x"3976812a",
          4342 => x"1770892a",
          4343 => x"a4180805",
          4344 => x"53765255",
          4345 => x"fb973f82",
          4346 => x"85ec0859",
          4347 => x"8285ec08",
          4348 => x"81d93874",
          4349 => x"83ff0616",
          4350 => x"b4058116",
          4351 => x"78810659",
          4352 => x"56547753",
          4353 => x"76802e8f",
          4354 => x"3877842b",
          4355 => x"9ff00674",
          4356 => x"338f0671",
          4357 => x"07515372",
          4358 => x"7434810b",
          4359 => x"83173474",
          4360 => x"892aa417",
          4361 => x"08055275",
          4362 => x"51fad23f",
          4363 => x"8285ec08",
          4364 => x"598285ec",
          4365 => x"08819438",
          4366 => x"7483ff06",
          4367 => x"16b40578",
          4368 => x"842a5454",
          4369 => x"768f3877",
          4370 => x"882a7433",
          4371 => x"81f00671",
          4372 => x"8f060751",
          4373 => x"53727434",
          4374 => x"80ec3976",
          4375 => x"882aa417",
          4376 => x"08055275",
          4377 => x"51fa963f",
          4378 => x"8285ec08",
          4379 => x"598285ec",
          4380 => x"0880d838",
          4381 => x"7783ffff",
          4382 => x"06527610",
          4383 => x"83fe0676",
          4384 => x"05b40551",
          4385 => x"f79d3fbe",
          4386 => x"3976872a",
          4387 => x"a4170805",
          4388 => x"527551f9",
          4389 => x"e83f8285",
          4390 => x"ec085982",
          4391 => x"85ec08ab",
          4392 => x"3877f00a",
          4393 => x"0677822b",
          4394 => x"83fc0670",
          4395 => x"18b40570",
          4396 => x"54515454",
          4397 => x"f6c23f82",
          4398 => x"85ec088f",
          4399 => x"0a067407",
          4400 => x"527251f6",
          4401 => x"fc3f810b",
          4402 => x"83173478",
          4403 => x"8285ec0c",
          4404 => x"8a3d0d04",
          4405 => x"f83d0d7a",
          4406 => x"7c7e7208",
          4407 => x"59565659",
          4408 => x"817527a4",
          4409 => x"38749817",
          4410 => x"08279d38",
          4411 => x"73802eaa",
          4412 => x"38ff5373",
          4413 => x"527551fd",
          4414 => x"a43f8285",
          4415 => x"ec085482",
          4416 => x"85ec0880",
          4417 => x"f2389339",
          4418 => x"825480eb",
          4419 => x"39815480",
          4420 => x"e6398285",
          4421 => x"ec085480",
          4422 => x"de397452",
          4423 => x"7851fb84",
          4424 => x"3f8285ec",
          4425 => x"08588285",
          4426 => x"ec08802e",
          4427 => x"80c73882",
          4428 => x"85ec0881",
          4429 => x"2ed23882",
          4430 => x"85ec08ff",
          4431 => x"2ecf3880",
          4432 => x"53745275",
          4433 => x"51fcd63f",
          4434 => x"8285ec08",
          4435 => x"c5389816",
          4436 => x"08fe1190",
          4437 => x"18085755",
          4438 => x"57747427",
          4439 => x"90388115",
          4440 => x"90170c84",
          4441 => x"16338107",
          4442 => x"54738417",
          4443 => x"34775576",
          4444 => x"7826ffa6",
          4445 => x"38805473",
          4446 => x"8285ec0c",
          4447 => x"8a3d0d04",
          4448 => x"f63d0d7c",
          4449 => x"7e710859",
          4450 => x"5b5b7995",
          4451 => x"388c1708",
          4452 => x"5877802e",
          4453 => x"88389817",
          4454 => x"087826b2",
          4455 => x"388158ae",
          4456 => x"3979527a",
          4457 => x"51f9fd3f",
          4458 => x"81557482",
          4459 => x"85ec0827",
          4460 => x"82e63882",
          4461 => x"85ec0855",
          4462 => x"8285ec08",
          4463 => x"ff2e82d8",
          4464 => x"38981708",
          4465 => x"8285ec08",
          4466 => x"2682cd38",
          4467 => x"79589017",
          4468 => x"08705654",
          4469 => x"73802e82",
          4470 => x"bf38777a",
          4471 => x"2e098106",
          4472 => x"80e43881",
          4473 => x"1a569817",
          4474 => x"08762683",
          4475 => x"38825675",
          4476 => x"527a51f9",
          4477 => x"af3f8059",
          4478 => x"8285ec08",
          4479 => x"812e0981",
          4480 => x"06863882",
          4481 => x"85ec0859",
          4482 => x"8285ec08",
          4483 => x"09700981",
          4484 => x"05707207",
          4485 => x"8025707c",
          4486 => x"078285ec",
          4487 => x"08545151",
          4488 => x"55557381",
          4489 => x"f3388285",
          4490 => x"ec08802e",
          4491 => x"95388c17",
          4492 => x"08548174",
          4493 => x"27903873",
          4494 => x"98180827",
          4495 => x"89387358",
          4496 => x"85397580",
          4497 => x"dd387756",
          4498 => x"81165698",
          4499 => x"17087626",
          4500 => x"89388256",
          4501 => x"75782681",
          4502 => x"b0387552",
          4503 => x"7a51f8c4",
          4504 => x"3f8285ec",
          4505 => x"08802eba",
          4506 => x"38805982",
          4507 => x"85ec0881",
          4508 => x"2e098106",
          4509 => x"86388285",
          4510 => x"ec085982",
          4511 => x"85ec0809",
          4512 => x"70098105",
          4513 => x"70720780",
          4514 => x"25707c07",
          4515 => x"51515555",
          4516 => x"7380fa38",
          4517 => x"75782e09",
          4518 => x"8106ffac",
          4519 => x"38735580",
          4520 => x"f739ff53",
          4521 => x"75527651",
          4522 => x"f9f33f82",
          4523 => x"85ec0882",
          4524 => x"85ec0809",
          4525 => x"81057082",
          4526 => x"85ec0807",
          4527 => x"80255155",
          4528 => x"5579802e",
          4529 => x"94387380",
          4530 => x"2e8f3875",
          4531 => x"53795276",
          4532 => x"51f9ca3f",
          4533 => x"8285ec08",
          4534 => x"5574a538",
          4535 => x"758c180c",
          4536 => x"981708fe",
          4537 => x"05901808",
          4538 => x"56547474",
          4539 => x"268638ff",
          4540 => x"1590180c",
          4541 => x"84173381",
          4542 => x"07547384",
          4543 => x"18349739",
          4544 => x"ff567481",
          4545 => x"2e90388c",
          4546 => x"3980558c",
          4547 => x"398285ec",
          4548 => x"08558539",
          4549 => x"81567555",
          4550 => x"748285ec",
          4551 => x"0c8c3d0d",
          4552 => x"04f83d0d",
          4553 => x"7a705255",
          4554 => x"f3e33f82",
          4555 => x"85ec0858",
          4556 => x"81568285",
          4557 => x"ec0880da",
          4558 => x"387b5274",
          4559 => x"51f6b43f",
          4560 => x"8285ec08",
          4561 => x"8285ec08",
          4562 => x"b0170c59",
          4563 => x"84805377",
          4564 => x"52b41570",
          4565 => x"5257f2bb",
          4566 => x"3f775684",
          4567 => x"39811656",
          4568 => x"8a152258",
          4569 => x"75782797",
          4570 => x"38815475",
          4571 => x"19537652",
          4572 => x"81153351",
          4573 => x"eddc3f82",
          4574 => x"85ec0880",
          4575 => x"2edf388a",
          4576 => x"15227632",
          4577 => x"70098105",
          4578 => x"70720770",
          4579 => x"9f2a5351",
          4580 => x"56567582",
          4581 => x"85ec0c8a",
          4582 => x"3d0d04f8",
          4583 => x"3d0d7a7c",
          4584 => x"71085856",
          4585 => x"5774f080",
          4586 => x"0a2680f1",
          4587 => x"38749f06",
          4588 => x"537280e9",
          4589 => x"38749018",
          4590 => x"0c881708",
          4591 => x"5473aa38",
          4592 => x"75335382",
          4593 => x"73278838",
          4594 => x"a8160854",
          4595 => x"739b3874",
          4596 => x"852a5382",
          4597 => x"0b881722",
          4598 => x"5a587279",
          4599 => x"2780fe38",
          4600 => x"a8160898",
          4601 => x"180c80cd",
          4602 => x"398a1622",
          4603 => x"70892b54",
          4604 => x"58727526",
          4605 => x"b2387352",
          4606 => x"7651f5a8",
          4607 => x"3f8285ec",
          4608 => x"08548285",
          4609 => x"ec08ff2e",
          4610 => x"bd38810b",
          4611 => x"8285ec08",
          4612 => x"278b3898",
          4613 => x"16088285",
          4614 => x"ec082685",
          4615 => x"388258bd",
          4616 => x"39747331",
          4617 => x"55cb3973",
          4618 => x"527551f4",
          4619 => x"c63f8285",
          4620 => x"ec089818",
          4621 => x"0c739418",
          4622 => x"0c981708",
          4623 => x"53825872",
          4624 => x"802e9a38",
          4625 => x"85398158",
          4626 => x"94397489",
          4627 => x"2a139818",
          4628 => x"0c7483ff",
          4629 => x"0616b405",
          4630 => x"9c180c80",
          4631 => x"58778285",
          4632 => x"ec0c8a3d",
          4633 => x"0d04f83d",
          4634 => x"0d7a7008",
          4635 => x"901208a0",
          4636 => x"05595754",
          4637 => x"f0800a77",
          4638 => x"27863880",
          4639 => x"0b98150c",
          4640 => x"98140853",
          4641 => x"84557280",
          4642 => x"2e81cb38",
          4643 => x"7683ff06",
          4644 => x"587781b5",
          4645 => x"38811398",
          4646 => x"150c9414",
          4647 => x"08557492",
          4648 => x"3876852a",
          4649 => x"88172256",
          4650 => x"53747326",
          4651 => x"819b3880",
          4652 => x"c0398a16",
          4653 => x"22ff0577",
          4654 => x"892a0653",
          4655 => x"72818a38",
          4656 => x"74527351",
          4657 => x"f3de3f82",
          4658 => x"85ec0853",
          4659 => x"8255810b",
          4660 => x"8285ec08",
          4661 => x"2780ff38",
          4662 => x"81558285",
          4663 => x"ec08ff2e",
          4664 => x"80f43898",
          4665 => x"16088285",
          4666 => x"ec082680",
          4667 => x"ca387b8a",
          4668 => x"38779815",
          4669 => x"0c845580",
          4670 => x"dd399414",
          4671 => x"08527351",
          4672 => x"f8fe3f82",
          4673 => x"85ec0853",
          4674 => x"87558285",
          4675 => x"ec08802e",
          4676 => x"80c43882",
          4677 => x"558285ec",
          4678 => x"08812eba",
          4679 => x"38815582",
          4680 => x"85ec08ff",
          4681 => x"2eb03882",
          4682 => x"85ec0852",
          4683 => x"7551fbf1",
          4684 => x"3f8285ec",
          4685 => x"08a03872",
          4686 => x"94150c72",
          4687 => x"527551f2",
          4688 => x"b23f8285",
          4689 => x"ec089815",
          4690 => x"0c769015",
          4691 => x"0c7716b4",
          4692 => x"059c150c",
          4693 => x"80557482",
          4694 => x"85ec0c8a",
          4695 => x"3d0d04f7",
          4696 => x"3d0d7b7d",
          4697 => x"71085b5b",
          4698 => x"57805276",
          4699 => x"51fcac3f",
          4700 => x"8285ec08",
          4701 => x"548285ec",
          4702 => x"0880ec38",
          4703 => x"8285ec08",
          4704 => x"56981708",
          4705 => x"527851ef",
          4706 => x"f43f8285",
          4707 => x"ec085482",
          4708 => x"85ec0880",
          4709 => x"d2388285",
          4710 => x"ec089c18",
          4711 => x"08703351",
          4712 => x"54587281",
          4713 => x"e52e0981",
          4714 => x"06833881",
          4715 => x"588285ec",
          4716 => x"08557283",
          4717 => x"38815577",
          4718 => x"75075372",
          4719 => x"802e8e38",
          4720 => x"81165675",
          4721 => x"7a2e0981",
          4722 => x"068838a5",
          4723 => x"398285ec",
          4724 => x"08568152",
          4725 => x"7651fd8e",
          4726 => x"3f8285ec",
          4727 => x"08548285",
          4728 => x"ec08802e",
          4729 => x"ff9b3873",
          4730 => x"842e0981",
          4731 => x"06833887",
          4732 => x"54738285",
          4733 => x"ec0c8b3d",
          4734 => x"0d04fd3d",
          4735 => x"0d769a11",
          4736 => x"5254ebdd",
          4737 => x"3f8285ec",
          4738 => x"0883ffff",
          4739 => x"06767033",
          4740 => x"51535371",
          4741 => x"832e0981",
          4742 => x"06903894",
          4743 => x"1451ebc1",
          4744 => x"3f8285ec",
          4745 => x"08902b73",
          4746 => x"07537282",
          4747 => x"85ec0c85",
          4748 => x"3d0d04fc",
          4749 => x"3d0d7779",
          4750 => x"7083ffff",
          4751 => x"06549a12",
          4752 => x"535555eb",
          4753 => x"de3f7670",
          4754 => x"33515372",
          4755 => x"832e0981",
          4756 => x"068b3873",
          4757 => x"902a5294",
          4758 => x"1551ebc7",
          4759 => x"3f863d0d",
          4760 => x"04f73d0d",
          4761 => x"7b7d5b55",
          4762 => x"8475085a",
          4763 => x"58981508",
          4764 => x"802e818a",
          4765 => x"38981508",
          4766 => x"527851ee",
          4767 => x"803f8285",
          4768 => x"ec085882",
          4769 => x"85ec0880",
          4770 => x"f5389c15",
          4771 => x"08703355",
          4772 => x"53738638",
          4773 => x"845880e6",
          4774 => x"398b1333",
          4775 => x"70bf0670",
          4776 => x"81ff0658",
          4777 => x"51537286",
          4778 => x"16348285",
          4779 => x"ec085373",
          4780 => x"81e52e83",
          4781 => x"38815373",
          4782 => x"ae2ea938",
          4783 => x"81707406",
          4784 => x"54577280",
          4785 => x"2e9e3875",
          4786 => x"8f2e9938",
          4787 => x"8285ec08",
          4788 => x"76df0654",
          4789 => x"5472882e",
          4790 => x"09810683",
          4791 => x"38765473",
          4792 => x"7a2ea038",
          4793 => x"80527451",
          4794 => x"fafc3f82",
          4795 => x"85ec0858",
          4796 => x"8285ec08",
          4797 => x"89389815",
          4798 => x"08fefa38",
          4799 => x"8639800b",
          4800 => x"98160c77",
          4801 => x"8285ec0c",
          4802 => x"8b3d0d04",
          4803 => x"fb3d0d77",
          4804 => x"70085754",
          4805 => x"81527351",
          4806 => x"fcc53f82",
          4807 => x"85ec0855",
          4808 => x"8285ec08",
          4809 => x"b4389814",
          4810 => x"08527551",
          4811 => x"eccf3f82",
          4812 => x"85ec0855",
          4813 => x"8285ec08",
          4814 => x"a038a053",
          4815 => x"8285ec08",
          4816 => x"529c1408",
          4817 => x"51eacc3f",
          4818 => x"8b53a014",
          4819 => x"529c1408",
          4820 => x"51ea9d3f",
          4821 => x"810b8317",
          4822 => x"34748285",
          4823 => x"ec0c873d",
          4824 => x"0d04fd3d",
          4825 => x"0d757008",
          4826 => x"98120854",
          4827 => x"70535553",
          4828 => x"ec8b3f82",
          4829 => x"85ec088d",
          4830 => x"389c1308",
          4831 => x"53e57334",
          4832 => x"810b8315",
          4833 => x"34853d0d",
          4834 => x"04fa3d0d",
          4835 => x"787a5757",
          4836 => x"800b8917",
          4837 => x"34981708",
          4838 => x"802e8182",
          4839 => x"38807089",
          4840 => x"18555555",
          4841 => x"9c170814",
          4842 => x"70338116",
          4843 => x"56515271",
          4844 => x"a02ea838",
          4845 => x"71852e09",
          4846 => x"81068438",
          4847 => x"81e55273",
          4848 => x"892e0981",
          4849 => x"068b38ae",
          4850 => x"73708105",
          4851 => x"55348115",
          4852 => x"55717370",
          4853 => x"81055534",
          4854 => x"8115558a",
          4855 => x"7427c538",
          4856 => x"75158805",
          4857 => x"52800b81",
          4858 => x"13349c17",
          4859 => x"08528b12",
          4860 => x"33881734",
          4861 => x"9c17089c",
          4862 => x"115252e7",
          4863 => x"fb3f8285",
          4864 => x"ec08760c",
          4865 => x"961251e7",
          4866 => x"d83f8285",
          4867 => x"ec088617",
          4868 => x"23981251",
          4869 => x"e7cb3f82",
          4870 => x"85ec0884",
          4871 => x"1723883d",
          4872 => x"0d04f33d",
          4873 => x"0d7f7008",
          4874 => x"5e5b8061",
          4875 => x"70335155",
          4876 => x"5573af2e",
          4877 => x"83388155",
          4878 => x"7380dc2e",
          4879 => x"91387480",
          4880 => x"2e8c3894",
          4881 => x"1d08881c",
          4882 => x"0cac3981",
          4883 => x"15418061",
          4884 => x"70335656",
          4885 => x"5673af2e",
          4886 => x"09810683",
          4887 => x"38815673",
          4888 => x"80dc3270",
          4889 => x"09810570",
          4890 => x"80257807",
          4891 => x"51515473",
          4892 => x"da387388",
          4893 => x"1c0c6070",
          4894 => x"33515473",
          4895 => x"9f269638",
          4896 => x"ff800bab",
          4897 => x"1c348052",
          4898 => x"7a51f68f",
          4899 => x"3f8285ec",
          4900 => x"085585a6",
          4901 => x"39913d61",
          4902 => x"a01d5c5a",
          4903 => x"5e8b53a0",
          4904 => x"527951e7",
          4905 => x"ee3f8070",
          4906 => x"59578879",
          4907 => x"33555c73",
          4908 => x"ae2e0981",
          4909 => x"0680d838",
          4910 => x"78187033",
          4911 => x"811a71ae",
          4912 => x"32700981",
          4913 => x"05709f2a",
          4914 => x"73822607",
          4915 => x"5151535a",
          4916 => x"5754738c",
          4917 => x"38791754",
          4918 => x"75743481",
          4919 => x"1757d939",
          4920 => x"75af3270",
          4921 => x"09810570",
          4922 => x"9f2a5151",
          4923 => x"547580dc",
          4924 => x"2e8c3873",
          4925 => x"802e8738",
          4926 => x"75a02682",
          4927 => x"c7387719",
          4928 => x"7e0ca454",
          4929 => x"a0762782",
          4930 => x"c738a054",
          4931 => x"82c23978",
          4932 => x"18703381",
          4933 => x"1a5a5754",
          4934 => x"a0762782",
          4935 => x"863875af",
          4936 => x"32700981",
          4937 => x"057780dc",
          4938 => x"32700981",
          4939 => x"05728025",
          4940 => x"71802507",
          4941 => x"51515651",
          4942 => x"5573802e",
          4943 => x"ae388439",
          4944 => x"81185880",
          4945 => x"781a7033",
          4946 => x"51555573",
          4947 => x"af2e0981",
          4948 => x"06833881",
          4949 => x"557380dc",
          4950 => x"32700981",
          4951 => x"05708025",
          4952 => x"77075151",
          4953 => x"5473d938",
          4954 => x"81b93975",
          4955 => x"ae2e0981",
          4956 => x"06833881",
          4957 => x"54767c27",
          4958 => x"74075473",
          4959 => x"802ea638",
          4960 => x"7b8b3270",
          4961 => x"09810577",
          4962 => x"ae327009",
          4963 => x"81057280",
          4964 => x"25719f2a",
          4965 => x"07535156",
          4966 => x"51557481",
          4967 => x"a7388857",
          4968 => x"8b5cfeeb",
          4969 => x"3975982b",
          4970 => x"54738025",
          4971 => x"8c387580",
          4972 => x"ff0681ff",
          4973 => x"b4113357",
          4974 => x"547551e6",
          4975 => x"c23f8285",
          4976 => x"ec08802e",
          4977 => x"b2387818",
          4978 => x"7033811a",
          4979 => x"71545a56",
          4980 => x"54e6b33f",
          4981 => x"8285ec08",
          4982 => x"802e80e8",
          4983 => x"38ff1c54",
          4984 => x"76742780",
          4985 => x"df387917",
          4986 => x"54757434",
          4987 => x"81177a11",
          4988 => x"55577474",
          4989 => x"34a73975",
          4990 => x"5281fed4",
          4991 => x"51e5df3f",
          4992 => x"8285ec08",
          4993 => x"bf38ff9f",
          4994 => x"16547399",
          4995 => x"268938e0",
          4996 => x"167081ff",
          4997 => x"06575479",
          4998 => x"17547574",
          4999 => x"34811757",
          5000 => x"fded3977",
          5001 => x"197e0c76",
          5002 => x"802e9938",
          5003 => x"79335473",
          5004 => x"81e52e09",
          5005 => x"81068438",
          5006 => x"857a3484",
          5007 => x"54a07627",
          5008 => x"8f388b39",
          5009 => x"865581f2",
          5010 => x"39845680",
          5011 => x"f3398054",
          5012 => x"738b1b34",
          5013 => x"807b0858",
          5014 => x"527a51f2",
          5015 => x"be3f8285",
          5016 => x"ec085682",
          5017 => x"85ec0880",
          5018 => x"d738981b",
          5019 => x"08527651",
          5020 => x"e68b3f82",
          5021 => x"85ec0856",
          5022 => x"8285ec08",
          5023 => x"80c2389c",
          5024 => x"1b087033",
          5025 => x"55557380",
          5026 => x"2effbe38",
          5027 => x"8b1533bf",
          5028 => x"06547386",
          5029 => x"1c348b15",
          5030 => x"3370832a",
          5031 => x"70810651",
          5032 => x"55587392",
          5033 => x"388b5379",
          5034 => x"527451e4",
          5035 => x"803f8285",
          5036 => x"ec08802e",
          5037 => x"8b387552",
          5038 => x"7a51f3aa",
          5039 => x"3fff9f39",
          5040 => x"75ab1c33",
          5041 => x"57557480",
          5042 => x"2ebb3874",
          5043 => x"842e0981",
          5044 => x"0680e738",
          5045 => x"75852a70",
          5046 => x"81067782",
          5047 => x"2a585154",
          5048 => x"73802e96",
          5049 => x"38758106",
          5050 => x"5473802e",
          5051 => x"fba738ff",
          5052 => x"800bab1c",
          5053 => x"34805580",
          5054 => x"c1397581",
          5055 => x"065473ba",
          5056 => x"388555b6",
          5057 => x"3975822a",
          5058 => x"70810651",
          5059 => x"5473ab38",
          5060 => x"861b3370",
          5061 => x"842a7081",
          5062 => x"06515555",
          5063 => x"73802ee1",
          5064 => x"38901b08",
          5065 => x"83ff061d",
          5066 => x"b405527c",
          5067 => x"51f5cb3f",
          5068 => x"8285ec08",
          5069 => x"881c0cfa",
          5070 => x"dc397482",
          5071 => x"85ec0c8f",
          5072 => x"3d0d04f6",
          5073 => x"3d0d7c5b",
          5074 => x"ff7b0870",
          5075 => x"71735559",
          5076 => x"5c555973",
          5077 => x"802e81cc",
          5078 => x"38757081",
          5079 => x"05573370",
          5080 => x"a0265252",
          5081 => x"71ba2e8d",
          5082 => x"3870ee38",
          5083 => x"71ba2e09",
          5084 => x"810681ab",
          5085 => x"387333d0",
          5086 => x"117081ff",
          5087 => x"06515253",
          5088 => x"70892691",
          5089 => x"38821473",
          5090 => x"81ff06d0",
          5091 => x"05565271",
          5092 => x"762e80fd",
          5093 => x"38800b81",
          5094 => x"ffa45955",
          5095 => x"77087a55",
          5096 => x"57767081",
          5097 => x"05583374",
          5098 => x"70810556",
          5099 => x"33ff9f12",
          5100 => x"53535370",
          5101 => x"99268938",
          5102 => x"e0137081",
          5103 => x"ff065451",
          5104 => x"ff9f1251",
          5105 => x"70992689",
          5106 => x"38e01270",
          5107 => x"81ff0653",
          5108 => x"51720981",
          5109 => x"05709f2a",
          5110 => x"51517272",
          5111 => x"2e098106",
          5112 => x"853870ff",
          5113 => x"bc387209",
          5114 => x"81057477",
          5115 => x"32700981",
          5116 => x"05707207",
          5117 => x"9f2a739f",
          5118 => x"2a075354",
          5119 => x"54517080",
          5120 => x"2e8f3881",
          5121 => x"15841959",
          5122 => x"55837525",
          5123 => x"ff8e388b",
          5124 => x"39748324",
          5125 => x"86387476",
          5126 => x"7c0c5978",
          5127 => x"51863982",
          5128 => x"9da43351",
          5129 => x"708285ec",
          5130 => x"0c8c3d0d",
          5131 => x"04fa3d0d",
          5132 => x"7856800b",
          5133 => x"831734ff",
          5134 => x"0bb0170c",
          5135 => x"79527551",
          5136 => x"e2bb3f84",
          5137 => x"558285ec",
          5138 => x"08818238",
          5139 => x"84b21651",
          5140 => x"df8f3f82",
          5141 => x"85ec0883",
          5142 => x"ffff0654",
          5143 => x"83557382",
          5144 => x"d4d52e09",
          5145 => x"810680e5",
          5146 => x"38800bb4",
          5147 => x"17335657",
          5148 => x"7481e92e",
          5149 => x"09810683",
          5150 => x"38815774",
          5151 => x"81eb3270",
          5152 => x"09810570",
          5153 => x"80257907",
          5154 => x"51515473",
          5155 => x"8a387481",
          5156 => x"e82e0981",
          5157 => x"06b53883",
          5158 => x"5381fee4",
          5159 => x"5280ea16",
          5160 => x"51e08a3f",
          5161 => x"8285ec08",
          5162 => x"558285ec",
          5163 => x"08802e9d",
          5164 => x"38855381",
          5165 => x"fee85281",
          5166 => x"861651df",
          5167 => x"f03f8285",
          5168 => x"ec085582",
          5169 => x"85ec0880",
          5170 => x"2e833882",
          5171 => x"55748285",
          5172 => x"ec0c883d",
          5173 => x"0d04f13d",
          5174 => x"0d620284",
          5175 => x"0580cf05",
          5176 => x"33585580",
          5177 => x"750c6151",
          5178 => x"fcd93f82",
          5179 => x"85ec0858",
          5180 => x"8b56800b",
          5181 => x"8285ec08",
          5182 => x"24878338",
          5183 => x"8285ec08",
          5184 => x"822b829d",
          5185 => x"90110855",
          5186 => x"538c5673",
          5187 => x"802e86ee",
          5188 => x"3873750c",
          5189 => x"7681fe06",
          5190 => x"74335457",
          5191 => x"72802eae",
          5192 => x"38811433",
          5193 => x"51d7a43f",
          5194 => x"8285ec08",
          5195 => x"81ff0670",
          5196 => x"81065455",
          5197 => x"72983876",
          5198 => x"802e86c0",
          5199 => x"3874822a",
          5200 => x"70810651",
          5201 => x"538a5672",
          5202 => x"86b43886",
          5203 => x"af398074",
          5204 => x"34778115",
          5205 => x"34815281",
          5206 => x"143351d7",
          5207 => x"8c3f8285",
          5208 => x"ec0881ff",
          5209 => x"06708106",
          5210 => x"54558356",
          5211 => x"72868f38",
          5212 => x"76802e8f",
          5213 => x"3874822a",
          5214 => x"70810651",
          5215 => x"538a5672",
          5216 => x"85fc3880",
          5217 => x"70537452",
          5218 => x"5cfda23f",
          5219 => x"8285ec08",
          5220 => x"81ff0657",
          5221 => x"76822e09",
          5222 => x"810680e2",
          5223 => x"388d3d74",
          5224 => x"56588356",
          5225 => x"83f61533",
          5226 => x"70585372",
          5227 => x"802e8d38",
          5228 => x"83fa1551",
          5229 => x"dcc23f82",
          5230 => x"85ec0857",
          5231 => x"76787084",
          5232 => x"055a0cff",
          5233 => x"16901656",
          5234 => x"56758025",
          5235 => x"d738800b",
          5236 => x"8e3d5456",
          5237 => x"72708405",
          5238 => x"54085c83",
          5239 => x"577b802e",
          5240 => x"95387b52",
          5241 => x"7351fcc5",
          5242 => x"3f8285ec",
          5243 => x"0881ff06",
          5244 => x"57817727",
          5245 => x"89388116",
          5246 => x"56837627",
          5247 => x"d7388156",
          5248 => x"76842e84",
          5249 => x"f9388d56",
          5250 => x"76812684",
          5251 => x"f138bf14",
          5252 => x"51dbce3f",
          5253 => x"8285ec08",
          5254 => x"83ffff06",
          5255 => x"53728480",
          5256 => x"2e098106",
          5257 => x"84d83880",
          5258 => x"ca1451db",
          5259 => x"b43f8285",
          5260 => x"ec0883ff",
          5261 => x"ff065877",
          5262 => x"8d3880d8",
          5263 => x"1451dbb8",
          5264 => x"3f8285ec",
          5265 => x"0858779c",
          5266 => x"150c80c4",
          5267 => x"14338215",
          5268 => x"3480c414",
          5269 => x"33ff1170",
          5270 => x"81ff0651",
          5271 => x"54558d56",
          5272 => x"72812684",
          5273 => x"99387481",
          5274 => x"ff065277",
          5275 => x"51fef89a",
          5276 => x"3f8285ec",
          5277 => x"0880c115",
          5278 => x"33545872",
          5279 => x"8a152372",
          5280 => x"802e8b38",
          5281 => x"ff137306",
          5282 => x"5372802e",
          5283 => x"86388d56",
          5284 => x"83ec3980",
          5285 => x"c51451da",
          5286 => x"c83f8285",
          5287 => x"ec085382",
          5288 => x"85ec0888",
          5289 => x"1523728f",
          5290 => x"06578d56",
          5291 => x"7683cf38",
          5292 => x"80c71451",
          5293 => x"daab3f82",
          5294 => x"85ec0883",
          5295 => x"ffff0655",
          5296 => x"748d3880",
          5297 => x"d41451da",
          5298 => x"af3f8285",
          5299 => x"ec085580",
          5300 => x"c21451da",
          5301 => x"8c3f8285",
          5302 => x"ec0883ff",
          5303 => x"ff065a8d",
          5304 => x"5679802e",
          5305 => x"83983888",
          5306 => x"1422781b",
          5307 => x"71842a05",
          5308 => x"5a5b7875",
          5309 => x"26838738",
          5310 => x"8a142252",
          5311 => x"74793151",
          5312 => x"fef8873f",
          5313 => x"8285ec08",
          5314 => x"538285ec",
          5315 => x"08802e82",
          5316 => x"ed388285",
          5317 => x"ec0880ff",
          5318 => x"fffff526",
          5319 => x"83388357",
          5320 => x"7283fff5",
          5321 => x"26833882",
          5322 => x"57729ff5",
          5323 => x"26853881",
          5324 => x"5789398d",
          5325 => x"5676802e",
          5326 => x"82c43882",
          5327 => x"13709816",
          5328 => x"0c7ca016",
          5329 => x"0c7a1d70",
          5330 => x"a4170c7a",
          5331 => x"1eac170c",
          5332 => x"54557683",
          5333 => x"2e098106",
          5334 => x"af3880de",
          5335 => x"1451d981",
          5336 => x"3f8285ec",
          5337 => x"0883ffff",
          5338 => x"06538d56",
          5339 => x"72828f38",
          5340 => x"7a828b38",
          5341 => x"80e01451",
          5342 => x"d8fe3f82",
          5343 => x"85ec08a8",
          5344 => x"150c7482",
          5345 => x"2b53a339",
          5346 => x"8d567a80",
          5347 => x"2e81ef38",
          5348 => x"7713a815",
          5349 => x"0c741553",
          5350 => x"76822e8e",
          5351 => x"38741075",
          5352 => x"11812a76",
          5353 => x"81061151",
          5354 => x"515383ff",
          5355 => x"13892a53",
          5356 => x"8d56729c",
          5357 => x"15082681",
          5358 => x"c538ff0b",
          5359 => x"90150cff",
          5360 => x"0b8c150c",
          5361 => x"ff800b84",
          5362 => x"15347683",
          5363 => x"2e098106",
          5364 => x"81923880",
          5365 => x"e41451d8",
          5366 => x"883f8285",
          5367 => x"ec0883ff",
          5368 => x"ff065372",
          5369 => x"812e0981",
          5370 => x"0680f938",
          5371 => x"811c5273",
          5372 => x"51db8a3f",
          5373 => x"8285ec08",
          5374 => x"80ea3882",
          5375 => x"85ec0884",
          5376 => x"153484b2",
          5377 => x"1451d7d9",
          5378 => x"3f8285ec",
          5379 => x"0883ffff",
          5380 => x"06537282",
          5381 => x"d4d52e09",
          5382 => x"810680c8",
          5383 => x"38b41451",
          5384 => x"d7d63f82",
          5385 => x"85ec0884",
          5386 => x"8b85a4d2",
          5387 => x"2e098106",
          5388 => x"b3388498",
          5389 => x"1451d7c0",
          5390 => x"3f8285ec",
          5391 => x"08868a85",
          5392 => x"e4f22e09",
          5393 => x"81069d38",
          5394 => x"849c1451",
          5395 => x"d7aa3f82",
          5396 => x"85ec0890",
          5397 => x"150c84a0",
          5398 => x"1451d79c",
          5399 => x"3f8285ec",
          5400 => x"088c150c",
          5401 => x"76743482",
          5402 => x"9da02281",
          5403 => x"05537282",
          5404 => x"9da02372",
          5405 => x"86152380",
          5406 => x"0b94150c",
          5407 => x"80567582",
          5408 => x"85ec0c91",
          5409 => x"3d0d04fb",
          5410 => x"3d0d7754",
          5411 => x"89557380",
          5412 => x"2eb93873",
          5413 => x"08537280",
          5414 => x"2eb13872",
          5415 => x"33527180",
          5416 => x"2ea93886",
          5417 => x"13228415",
          5418 => x"22575271",
          5419 => x"762e0981",
          5420 => x"06993881",
          5421 => x"133351d0",
          5422 => x"923f8285",
          5423 => x"ec088106",
          5424 => x"52718838",
          5425 => x"71740854",
          5426 => x"55833980",
          5427 => x"53787371",
          5428 => x"0c527482",
          5429 => x"85ec0c87",
          5430 => x"3d0d04fa",
          5431 => x"3d0d02ab",
          5432 => x"05337a58",
          5433 => x"893dfc05",
          5434 => x"5256f4d7",
          5435 => x"3f8b5480",
          5436 => x"0b8285ec",
          5437 => x"0824bc38",
          5438 => x"8285ec08",
          5439 => x"822b829d",
          5440 => x"90057008",
          5441 => x"55557380",
          5442 => x"2e843880",
          5443 => x"74347854",
          5444 => x"73802e84",
          5445 => x"38807434",
          5446 => x"78750c75",
          5447 => x"5475802e",
          5448 => x"92388053",
          5449 => x"893d7053",
          5450 => x"840551f7",
          5451 => x"a93f8285",
          5452 => x"ec085473",
          5453 => x"8285ec0c",
          5454 => x"883d0d04",
          5455 => x"eb3d0d67",
          5456 => x"02840580",
          5457 => x"e7053359",
          5458 => x"59895478",
          5459 => x"802e84ca",
          5460 => x"3877bf06",
          5461 => x"7054983d",
          5462 => x"d0055399",
          5463 => x"3d840552",
          5464 => x"58f6f33f",
          5465 => x"8285ec08",
          5466 => x"558285ec",
          5467 => x"0884a638",
          5468 => x"7a5c6852",
          5469 => x"8c3d7052",
          5470 => x"56eda73f",
          5471 => x"8285ec08",
          5472 => x"558285ec",
          5473 => x"08923802",
          5474 => x"80d70533",
          5475 => x"70982b55",
          5476 => x"57738025",
          5477 => x"83388655",
          5478 => x"779c0654",
          5479 => x"73802e81",
          5480 => x"ab387480",
          5481 => x"2e953874",
          5482 => x"842e0981",
          5483 => x"06aa3875",
          5484 => x"51ead93f",
          5485 => x"8285ec08",
          5486 => x"559e3902",
          5487 => x"b2053391",
          5488 => x"06547381",
          5489 => x"b8387782",
          5490 => x"2a708106",
          5491 => x"51547380",
          5492 => x"2e8e3888",
          5493 => x"5583be39",
          5494 => x"77880758",
          5495 => x"7483b638",
          5496 => x"77832a70",
          5497 => x"81065154",
          5498 => x"73802e81",
          5499 => x"af386252",
          5500 => x"7a51e886",
          5501 => x"3f8285ec",
          5502 => x"08568288",
          5503 => x"b20a5262",
          5504 => x"8e0551d4",
          5505 => x"bc3f6254",
          5506 => x"a00b8b15",
          5507 => x"34805362",
          5508 => x"527a51e8",
          5509 => x"9e3f8052",
          5510 => x"629c0551",
          5511 => x"d4a33f7a",
          5512 => x"54810b83",
          5513 => x"15347580",
          5514 => x"2e80f138",
          5515 => x"7ab01108",
          5516 => x"51548053",
          5517 => x"7552973d",
          5518 => x"d40551dd",
          5519 => x"973f8285",
          5520 => x"ec085582",
          5521 => x"85ec0882",
          5522 => x"cc38b739",
          5523 => x"7482c638",
          5524 => x"02b20533",
          5525 => x"70842a70",
          5526 => x"81065155",
          5527 => x"5673802e",
          5528 => x"86388455",
          5529 => x"82af3977",
          5530 => x"812a7081",
          5531 => x"06515473",
          5532 => x"802ea938",
          5533 => x"75810654",
          5534 => x"73802ea0",
          5535 => x"38875582",
          5536 => x"94397352",
          5537 => x"7a51d5f5",
          5538 => x"3f8285ec",
          5539 => x"087bff18",
          5540 => x"8c120c55",
          5541 => x"558285ec",
          5542 => x"0881fa38",
          5543 => x"77832a70",
          5544 => x"81065154",
          5545 => x"73802e86",
          5546 => x"387780c0",
          5547 => x"07587ab0",
          5548 => x"1108a01b",
          5549 => x"0c63a41b",
          5550 => x"0c635370",
          5551 => x"5257e6ba",
          5552 => x"3f8285ec",
          5553 => x"088285ec",
          5554 => x"08881b0c",
          5555 => x"639c0552",
          5556 => x"5ad2a53f",
          5557 => x"8285ec08",
          5558 => x"8285ec08",
          5559 => x"8c1b0c77",
          5560 => x"7a0c5686",
          5561 => x"1722841a",
          5562 => x"2377901a",
          5563 => x"34800b91",
          5564 => x"1a34800b",
          5565 => x"9c1a0c80",
          5566 => x"0b941a0c",
          5567 => x"77852a70",
          5568 => x"81065154",
          5569 => x"73802e81",
          5570 => x"8f388285",
          5571 => x"ec08802e",
          5572 => x"81863882",
          5573 => x"85ec0894",
          5574 => x"1a0c8a17",
          5575 => x"2270892b",
          5576 => x"7b525957",
          5577 => x"a8397652",
          5578 => x"7851d6f8",
          5579 => x"3f8285ec",
          5580 => x"08578285",
          5581 => x"ec088126",
          5582 => x"83388255",
          5583 => x"8285ec08",
          5584 => x"ff2e0981",
          5585 => x"06833879",
          5586 => x"55757831",
          5587 => x"56740981",
          5588 => x"05707607",
          5589 => x"80255154",
          5590 => x"7776278a",
          5591 => x"38817075",
          5592 => x"06555a73",
          5593 => x"c1387698",
          5594 => x"1a0c74a9",
          5595 => x"387583ff",
          5596 => x"06547380",
          5597 => x"2ea23876",
          5598 => x"527a51d5",
          5599 => x"f63f8285",
          5600 => x"ec088538",
          5601 => x"82558e39",
          5602 => x"75892a82",
          5603 => x"85ec0805",
          5604 => x"9c1a0c84",
          5605 => x"3980790c",
          5606 => x"74547382",
          5607 => x"85ec0c97",
          5608 => x"3d0d04f2",
          5609 => x"3d0d6063",
          5610 => x"65644040",
          5611 => x"5d59807e",
          5612 => x"0c903dfc",
          5613 => x"05527851",
          5614 => x"f9cd3f82",
          5615 => x"85ec0855",
          5616 => x"8285ec08",
          5617 => x"8a389119",
          5618 => x"33557480",
          5619 => x"2e863874",
          5620 => x"5682c439",
          5621 => x"90193381",
          5622 => x"06558756",
          5623 => x"74802e82",
          5624 => x"b6389539",
          5625 => x"820b911a",
          5626 => x"34825682",
          5627 => x"aa39810b",
          5628 => x"911a3481",
          5629 => x"5682a039",
          5630 => x"8c190894",
          5631 => x"1a083155",
          5632 => x"747c2783",
          5633 => x"38745c7b",
          5634 => x"802e8289",
          5635 => x"38941908",
          5636 => x"7083ff06",
          5637 => x"56567481",
          5638 => x"b2387e8a",
          5639 => x"1122ff05",
          5640 => x"77892a06",
          5641 => x"5b5579a8",
          5642 => x"38758738",
          5643 => x"88190855",
          5644 => x"8f399819",
          5645 => x"08527851",
          5646 => x"d4ea3f82",
          5647 => x"85ec0855",
          5648 => x"817527ff",
          5649 => x"9f3874ff",
          5650 => x"2effa338",
          5651 => x"74981a0c",
          5652 => x"98190852",
          5653 => x"7e51d49b",
          5654 => x"3f8285ec",
          5655 => x"08802eff",
          5656 => x"83388285",
          5657 => x"ec081a7c",
          5658 => x"892a5957",
          5659 => x"77802e80",
          5660 => x"d638771a",
          5661 => x"7f8a1122",
          5662 => x"585c5575",
          5663 => x"75278538",
          5664 => x"757a3158",
          5665 => x"77547653",
          5666 => x"7c52811b",
          5667 => x"3351c9d8",
          5668 => x"3f8285ec",
          5669 => x"08fed738",
          5670 => x"7e831133",
          5671 => x"56567480",
          5672 => x"2e9f38b0",
          5673 => x"16087731",
          5674 => x"55747827",
          5675 => x"94388480",
          5676 => x"53b41652",
          5677 => x"b0160877",
          5678 => x"31892b7d",
          5679 => x"0551cfb0",
          5680 => x"3f77892b",
          5681 => x"56b93976",
          5682 => x"9c1a0c94",
          5683 => x"190883ff",
          5684 => x"06848071",
          5685 => x"3157557b",
          5686 => x"76278338",
          5687 => x"7b569c19",
          5688 => x"08527e51",
          5689 => x"d1973f82",
          5690 => x"85ec08fe",
          5691 => x"81387553",
          5692 => x"94190883",
          5693 => x"ff061fb4",
          5694 => x"05527c51",
          5695 => x"cef23f7b",
          5696 => x"76317e08",
          5697 => x"177f0c76",
          5698 => x"1e941b08",
          5699 => x"18941c0c",
          5700 => x"5e5cfdf3",
          5701 => x"39805675",
          5702 => x"8285ec0c",
          5703 => x"903d0d04",
          5704 => x"f23d0d60",
          5705 => x"63656440",
          5706 => x"405d5880",
          5707 => x"7e0c903d",
          5708 => x"fc055277",
          5709 => x"51f6d03f",
          5710 => x"8285ec08",
          5711 => x"558285ec",
          5712 => x"088a3891",
          5713 => x"18335574",
          5714 => x"802e8638",
          5715 => x"745683b8",
          5716 => x"39901833",
          5717 => x"70812a70",
          5718 => x"81065156",
          5719 => x"56875674",
          5720 => x"802e83a4",
          5721 => x"38953982",
          5722 => x"0b911934",
          5723 => x"82568398",
          5724 => x"39810b91",
          5725 => x"19348156",
          5726 => x"838e3994",
          5727 => x"18087c11",
          5728 => x"56567476",
          5729 => x"27843875",
          5730 => x"095c7b80",
          5731 => x"2e82ec38",
          5732 => x"94180870",
          5733 => x"83ff0656",
          5734 => x"567481fd",
          5735 => x"387e8a11",
          5736 => x"22ff0577",
          5737 => x"892a065c",
          5738 => x"557abf38",
          5739 => x"758c3888",
          5740 => x"18085574",
          5741 => x"9c387a52",
          5742 => x"85399818",
          5743 => x"08527751",
          5744 => x"d7be3f82",
          5745 => x"85ec0855",
          5746 => x"8285ec08",
          5747 => x"802e82ab",
          5748 => x"3874812e",
          5749 => x"ff913874",
          5750 => x"ff2eff95",
          5751 => x"38749819",
          5752 => x"0c881808",
          5753 => x"85387488",
          5754 => x"190c7e55",
          5755 => x"b015089c",
          5756 => x"19082e09",
          5757 => x"81068d38",
          5758 => x"7451ce91",
          5759 => x"3f8285ec",
          5760 => x"08feee38",
          5761 => x"98180852",
          5762 => x"7e51d0e7",
          5763 => x"3f8285ec",
          5764 => x"08802efe",
          5765 => x"d2388285",
          5766 => x"ec081b7c",
          5767 => x"892a5a57",
          5768 => x"78802e80",
          5769 => x"d538781b",
          5770 => x"7f8a1122",
          5771 => x"585b5575",
          5772 => x"75278538",
          5773 => x"757b3159",
          5774 => x"78547653",
          5775 => x"7c52811a",
          5776 => x"3351c88e",
          5777 => x"3f8285ec",
          5778 => x"08fea638",
          5779 => x"7eb01108",
          5780 => x"78315656",
          5781 => x"7479279b",
          5782 => x"38848053",
          5783 => x"b0160877",
          5784 => x"31892b7d",
          5785 => x"0552b416",
          5786 => x"51cc853f",
          5787 => x"7e55800b",
          5788 => x"83163478",
          5789 => x"892b5680",
          5790 => x"db398c18",
          5791 => x"08941908",
          5792 => x"2693387e",
          5793 => x"51cd863f",
          5794 => x"8285ec08",
          5795 => x"fde3387e",
          5796 => x"77b0120c",
          5797 => x"55769c19",
          5798 => x"0c941808",
          5799 => x"83ff0684",
          5800 => x"80713157",
          5801 => x"557b7627",
          5802 => x"83387b56",
          5803 => x"9c180852",
          5804 => x"7e51cdc9",
          5805 => x"3f8285ec",
          5806 => x"08fdb638",
          5807 => x"75537c52",
          5808 => x"94180883",
          5809 => x"ff061fb4",
          5810 => x"0551cba4",
          5811 => x"3f7e5581",
          5812 => x"0b831634",
          5813 => x"7b76317e",
          5814 => x"08177f0c",
          5815 => x"761e941a",
          5816 => x"08187094",
          5817 => x"1c0c8c1b",
          5818 => x"0858585e",
          5819 => x"5c747627",
          5820 => x"83387555",
          5821 => x"748c190c",
          5822 => x"fd903990",
          5823 => x"183380c0",
          5824 => x"07557490",
          5825 => x"19348056",
          5826 => x"758285ec",
          5827 => x"0c903d0d",
          5828 => x"04f83d0d",
          5829 => x"7a8b3dfc",
          5830 => x"05537052",
          5831 => x"56f2e83f",
          5832 => x"8285ec08",
          5833 => x"578285ec",
          5834 => x"0880fb38",
          5835 => x"90163370",
          5836 => x"862a7081",
          5837 => x"06515555",
          5838 => x"73802e80",
          5839 => x"e938a016",
          5840 => x"08527851",
          5841 => x"ccb73f82",
          5842 => x"85ec0857",
          5843 => x"8285ec08",
          5844 => x"80d438a4",
          5845 => x"16088b11",
          5846 => x"33a00755",
          5847 => x"55738b16",
          5848 => x"34881608",
          5849 => x"53745275",
          5850 => x"0851ddc7",
          5851 => x"3f8c1608",
          5852 => x"529c1551",
          5853 => x"c9cb3f82",
          5854 => x"88b20a52",
          5855 => x"961551c9",
          5856 => x"c03f7652",
          5857 => x"921551c9",
          5858 => x"9a3f7854",
          5859 => x"810b8315",
          5860 => x"347851cc",
          5861 => x"af3f8285",
          5862 => x"ec089017",
          5863 => x"3381bf06",
          5864 => x"55577390",
          5865 => x"17347682",
          5866 => x"85ec0c8a",
          5867 => x"3d0d04fc",
          5868 => x"3d0d7670",
          5869 => x"5254fed9",
          5870 => x"3f8285ec",
          5871 => x"08538285",
          5872 => x"ec089c38",
          5873 => x"863dfc05",
          5874 => x"527351f1",
          5875 => x"ba3f8285",
          5876 => x"ec085382",
          5877 => x"85ec0887",
          5878 => x"388285ec",
          5879 => x"08740c72",
          5880 => x"8285ec0c",
          5881 => x"863d0d04",
          5882 => x"ff3d0d84",
          5883 => x"3d51e6d3",
          5884 => x"3f8b5280",
          5885 => x"0b8285ec",
          5886 => x"08248b38",
          5887 => x"8285ec08",
          5888 => x"829da434",
          5889 => x"80527182",
          5890 => x"85ec0c83",
          5891 => x"3d0d04ef",
          5892 => x"3d0d8053",
          5893 => x"933dd005",
          5894 => x"52943d51",
          5895 => x"e9b83f82",
          5896 => x"85ec0855",
          5897 => x"8285ec08",
          5898 => x"80e03876",
          5899 => x"58635293",
          5900 => x"3dd40551",
          5901 => x"dfec3f82",
          5902 => x"85ec0855",
          5903 => x"8285ec08",
          5904 => x"bc380280",
          5905 => x"c7053370",
          5906 => x"982b5556",
          5907 => x"73802589",
          5908 => x"38767a94",
          5909 => x"120c54b2",
          5910 => x"3902a205",
          5911 => x"3370842a",
          5912 => x"70810651",
          5913 => x"55567380",
          5914 => x"2e9e3876",
          5915 => x"7f537052",
          5916 => x"54db873f",
          5917 => x"8285ec08",
          5918 => x"94150c8e",
          5919 => x"398285ec",
          5920 => x"08842e09",
          5921 => x"81068338",
          5922 => x"85557482",
          5923 => x"85ec0c93",
          5924 => x"3d0d04e4",
          5925 => x"3d0d6f6f",
          5926 => x"5b5b807a",
          5927 => x"3480539e",
          5928 => x"3dffb805",
          5929 => x"529f3d51",
          5930 => x"e8ac3f82",
          5931 => x"85ec0857",
          5932 => x"8285ec08",
          5933 => x"82fb387b",
          5934 => x"437a7c94",
          5935 => x"11084755",
          5936 => x"58645473",
          5937 => x"802e81ed",
          5938 => x"38a05293",
          5939 => x"3d705255",
          5940 => x"d5c93f82",
          5941 => x"85ec0857",
          5942 => x"8285ec08",
          5943 => x"82d33868",
          5944 => x"527b51c9",
          5945 => x"983f8285",
          5946 => x"ec085782",
          5947 => x"85ec0882",
          5948 => x"c0386952",
          5949 => x"7b51da82",
          5950 => x"3f8285ec",
          5951 => x"08457652",
          5952 => x"7451d597",
          5953 => x"3f8285ec",
          5954 => x"08578285",
          5955 => x"ec0882a1",
          5956 => x"38805274",
          5957 => x"51daca3f",
          5958 => x"8285ec08",
          5959 => x"578285ec",
          5960 => x"08a43869",
          5961 => x"527b51d9",
          5962 => x"d13f7382",
          5963 => x"85ec082e",
          5964 => x"a6387652",
          5965 => x"7451d6ae",
          5966 => x"3f8285ec",
          5967 => x"08578285",
          5968 => x"ec08802e",
          5969 => x"cc387684",
          5970 => x"2e098106",
          5971 => x"86388257",
          5972 => x"81df3976",
          5973 => x"81db389e",
          5974 => x"3dffbc05",
          5975 => x"527451dc",
          5976 => x"a83f7690",
          5977 => x"3d781181",
          5978 => x"11335156",
          5979 => x"5a567380",
          5980 => x"2e913802",
          5981 => x"b9055581",
          5982 => x"16811670",
          5983 => x"33565656",
          5984 => x"73f53881",
          5985 => x"16547378",
          5986 => x"26818f38",
          5987 => x"75802e99",
          5988 => x"38781681",
          5989 => x"0555ff18",
          5990 => x"6f11ff18",
          5991 => x"ff185858",
          5992 => x"55587433",
          5993 => x"743475ee",
          5994 => x"38ff186f",
          5995 => x"115558af",
          5996 => x"7434fe8d",
          5997 => x"39777b2e",
          5998 => x"0981068a",
          5999 => x"38ff186f",
          6000 => x"115558af",
          6001 => x"7434800b",
          6002 => x"829da433",
          6003 => x"70822b81",
          6004 => x"ffa41108",
          6005 => x"7033525c",
          6006 => x"56565673",
          6007 => x"762e8d38",
          6008 => x"8116701a",
          6009 => x"70335155",
          6010 => x"5673f538",
          6011 => x"82165473",
          6012 => x"7826a738",
          6013 => x"80557476",
          6014 => x"27913874",
          6015 => x"19547333",
          6016 => x"7a708105",
          6017 => x"5c348115",
          6018 => x"55ec39ba",
          6019 => x"7a708105",
          6020 => x"5c3474ff",
          6021 => x"2e098106",
          6022 => x"85389157",
          6023 => x"94396e18",
          6024 => x"81195954",
          6025 => x"73337a70",
          6026 => x"81055c34",
          6027 => x"7a7826ee",
          6028 => x"38807a34",
          6029 => x"768285ec",
          6030 => x"0c9e3d0d",
          6031 => x"04f73d0d",
          6032 => x"7b7d8d3d",
          6033 => x"fc055471",
          6034 => x"535755ec",
          6035 => x"ba3f8285",
          6036 => x"ec085382",
          6037 => x"85ec0882",
          6038 => x"fc389115",
          6039 => x"33537282",
          6040 => x"f4388c15",
          6041 => x"08547376",
          6042 => x"27923890",
          6043 => x"15337081",
          6044 => x"2a708106",
          6045 => x"51545772",
          6046 => x"83387356",
          6047 => x"94150854",
          6048 => x"80709417",
          6049 => x"0c587578",
          6050 => x"2e829938",
          6051 => x"798a1122",
          6052 => x"70892b59",
          6053 => x"51537378",
          6054 => x"2eb93876",
          6055 => x"52ff1651",
          6056 => x"fee0e73f",
          6057 => x"8285ec08",
          6058 => x"ff157854",
          6059 => x"70535553",
          6060 => x"fee0d73f",
          6061 => x"8285ec08",
          6062 => x"73269838",
          6063 => x"76098105",
          6064 => x"70750670",
          6065 => x"94180c77",
          6066 => x"71319818",
          6067 => x"08575851",
          6068 => x"53b13988",
          6069 => x"15085473",
          6070 => x"a6387352",
          6071 => x"7451cda0",
          6072 => x"3f8285ec",
          6073 => x"08548285",
          6074 => x"ec08812e",
          6075 => x"819a3882",
          6076 => x"85ec08ff",
          6077 => x"2e819b38",
          6078 => x"8285ec08",
          6079 => x"88160c73",
          6080 => x"98160c73",
          6081 => x"802e819c",
          6082 => x"38767627",
          6083 => x"80dc3875",
          6084 => x"77319416",
          6085 => x"08189417",
          6086 => x"0c901633",
          6087 => x"70812a70",
          6088 => x"81065155",
          6089 => x"5a567280",
          6090 => x"2e9a3873",
          6091 => x"527451cc",
          6092 => x"cf3f8285",
          6093 => x"ec085482",
          6094 => x"85ec0894",
          6095 => x"388285ec",
          6096 => x"0856a739",
          6097 => x"73527451",
          6098 => x"c6da3f82",
          6099 => x"85ec0854",
          6100 => x"73ff2ebe",
          6101 => x"38817427",
          6102 => x"af387953",
          6103 => x"73981408",
          6104 => x"27a63873",
          6105 => x"98160cff",
          6106 => x"a0399415",
          6107 => x"08169416",
          6108 => x"0c7583ff",
          6109 => x"06537280",
          6110 => x"2eaa3873",
          6111 => x"527951c5",
          6112 => x"f23f8285",
          6113 => x"ec089438",
          6114 => x"820b9116",
          6115 => x"34825380",
          6116 => x"c439810b",
          6117 => x"91163481",
          6118 => x"53bb3975",
          6119 => x"892a8285",
          6120 => x"ec080558",
          6121 => x"94150854",
          6122 => x"8c150874",
          6123 => x"27903873",
          6124 => x"8c160c90",
          6125 => x"153380c0",
          6126 => x"07537290",
          6127 => x"16347383",
          6128 => x"ff065372",
          6129 => x"802e8c38",
          6130 => x"779c1608",
          6131 => x"2e853877",
          6132 => x"9c160c80",
          6133 => x"53728285",
          6134 => x"ec0c8b3d",
          6135 => x"0d04f93d",
          6136 => x"0d795689",
          6137 => x"5475802e",
          6138 => x"818a3880",
          6139 => x"53893dfc",
          6140 => x"05528a3d",
          6141 => x"840551e1",
          6142 => x"dd3f8285",
          6143 => x"ec085582",
          6144 => x"85ec0880",
          6145 => x"ea387776",
          6146 => x"0c7a5275",
          6147 => x"51d8933f",
          6148 => x"8285ec08",
          6149 => x"558285ec",
          6150 => x"0880c338",
          6151 => x"ab163370",
          6152 => x"982b5557",
          6153 => x"807424a2",
          6154 => x"38861633",
          6155 => x"70842a70",
          6156 => x"81065155",
          6157 => x"5773802e",
          6158 => x"ad389c16",
          6159 => x"08527751",
          6160 => x"d3b83f82",
          6161 => x"85ec0888",
          6162 => x"170c7754",
          6163 => x"86142284",
          6164 => x"17237452",
          6165 => x"7551cec3",
          6166 => x"3f8285ec",
          6167 => x"08557484",
          6168 => x"2e098106",
          6169 => x"85388555",
          6170 => x"86397480",
          6171 => x"2e843880",
          6172 => x"760c7454",
          6173 => x"738285ec",
          6174 => x"0c893d0d",
          6175 => x"04fc3d0d",
          6176 => x"76873dfc",
          6177 => x"05537052",
          6178 => x"53e7fc3f",
          6179 => x"8285ec08",
          6180 => x"87388285",
          6181 => x"ec08730c",
          6182 => x"863d0d04",
          6183 => x"fb3d0d77",
          6184 => x"79893dfc",
          6185 => x"05547153",
          6186 => x"5654e7db",
          6187 => x"3f8285ec",
          6188 => x"08538285",
          6189 => x"ec0880e1",
          6190 => x"38749338",
          6191 => x"8285ec08",
          6192 => x"527351cd",
          6193 => x"d63f8285",
          6194 => x"ec085380",
          6195 => x"cc398285",
          6196 => x"ec085273",
          6197 => x"51d38a3f",
          6198 => x"8285ec08",
          6199 => x"538285ec",
          6200 => x"08842e09",
          6201 => x"81068538",
          6202 => x"80538739",
          6203 => x"8285ec08",
          6204 => x"a8387452",
          6205 => x"7351d591",
          6206 => x"3f725273",
          6207 => x"51cee73f",
          6208 => x"8285ec08",
          6209 => x"84327009",
          6210 => x"81057072",
          6211 => x"079f2c70",
          6212 => x"8285ec08",
          6213 => x"06515154",
          6214 => x"54728285",
          6215 => x"ec0c873d",
          6216 => x"0d04ee3d",
          6217 => x"0d655780",
          6218 => x"53893d70",
          6219 => x"53963d52",
          6220 => x"56dfa33f",
          6221 => x"8285ec08",
          6222 => x"558285ec",
          6223 => x"08b23864",
          6224 => x"527551d5",
          6225 => x"dd3f8285",
          6226 => x"ec085582",
          6227 => x"85ec08a0",
          6228 => x"380280cb",
          6229 => x"05337098",
          6230 => x"2b555873",
          6231 => x"80258538",
          6232 => x"86558d39",
          6233 => x"76802e88",
          6234 => x"38765275",
          6235 => x"51d49a3f",
          6236 => x"748285ec",
          6237 => x"0c943d0d",
          6238 => x"04f03d0d",
          6239 => x"6365555c",
          6240 => x"8053923d",
          6241 => x"ec055293",
          6242 => x"3d51deca",
          6243 => x"3f8285ec",
          6244 => x"085b8285",
          6245 => x"ec088287",
          6246 => x"387c740c",
          6247 => x"73089811",
          6248 => x"08fe1190",
          6249 => x"13085956",
          6250 => x"58557574",
          6251 => x"26913875",
          6252 => x"7c0c81eb",
          6253 => x"39815b81",
          6254 => x"d339825b",
          6255 => x"81ce3982",
          6256 => x"85ec0875",
          6257 => x"33555973",
          6258 => x"812e0981",
          6259 => x"0680c138",
          6260 => x"82755f57",
          6261 => x"7652923d",
          6262 => x"f00551c1",
          6263 => x"c73f8285",
          6264 => x"ec08ff2e",
          6265 => x"d0388285",
          6266 => x"ec08812e",
          6267 => x"cd388285",
          6268 => x"ec080981",
          6269 => x"05708285",
          6270 => x"ec080780",
          6271 => x"257a0581",
          6272 => x"197f5359",
          6273 => x"5a549814",
          6274 => x"087726c8",
          6275 => x"3880fd39",
          6276 => x"a4150882",
          6277 => x"85ec0857",
          6278 => x"58759838",
          6279 => x"77528118",
          6280 => x"7d5258ff",
          6281 => x"bed73f82",
          6282 => x"85ec085b",
          6283 => x"8285ec08",
          6284 => x"80da387c",
          6285 => x"70337712",
          6286 => x"ff1a5d52",
          6287 => x"56547482",
          6288 => x"2e098106",
          6289 => x"a038b414",
          6290 => x"51ffbb95",
          6291 => x"3f8285ec",
          6292 => x"0883ffff",
          6293 => x"06700981",
          6294 => x"05708025",
          6295 => x"1b821959",
          6296 => x"5b51549d",
          6297 => x"39b41451",
          6298 => x"ffbb8d3f",
          6299 => x"8285ec08",
          6300 => x"f00a0670",
          6301 => x"09810570",
          6302 => x"80251b84",
          6303 => x"19595b51",
          6304 => x"547583ff",
          6305 => x"067a5856",
          6306 => x"79ff8e38",
          6307 => x"787c0c7c",
          6308 => x"7990120c",
          6309 => x"84113381",
          6310 => x"07565474",
          6311 => x"8415347a",
          6312 => x"8285ec0c",
          6313 => x"923d0d04",
          6314 => x"f93d0d79",
          6315 => x"8a3dfc05",
          6316 => x"53705257",
          6317 => x"e3d13f82",
          6318 => x"85ec0856",
          6319 => x"8285ec08",
          6320 => x"81a83891",
          6321 => x"17335675",
          6322 => x"81a03890",
          6323 => x"17337081",
          6324 => x"2a708106",
          6325 => x"51555587",
          6326 => x"5573802e",
          6327 => x"818e3894",
          6328 => x"17085473",
          6329 => x"8c180827",
          6330 => x"81803873",
          6331 => x"9b388285",
          6332 => x"ec085388",
          6333 => x"17085276",
          6334 => x"51c3d93f",
          6335 => x"8285ec08",
          6336 => x"7488190c",
          6337 => x"5680c939",
          6338 => x"98170852",
          6339 => x"7651ffbf",
          6340 => x"933f8285",
          6341 => x"ec08ff2e",
          6342 => x"09810683",
          6343 => x"38815682",
          6344 => x"85ec0881",
          6345 => x"2e098106",
          6346 => x"85388256",
          6347 => x"a33975a0",
          6348 => x"38775482",
          6349 => x"85ec0898",
          6350 => x"15082794",
          6351 => x"38981708",
          6352 => x"538285ec",
          6353 => x"08527651",
          6354 => x"c38a3f82",
          6355 => x"85ec0856",
          6356 => x"9417088c",
          6357 => x"180c9017",
          6358 => x"3380c007",
          6359 => x"54739018",
          6360 => x"3475802e",
          6361 => x"85387591",
          6362 => x"18347555",
          6363 => x"748285ec",
          6364 => x"0c893d0d",
          6365 => x"04e23d0d",
          6366 => x"8253a03d",
          6367 => x"ffa40552",
          6368 => x"a13d51da",
          6369 => x"d13f8285",
          6370 => x"ec085582",
          6371 => x"85ec0881",
          6372 => x"f7387845",
          6373 => x"a13d0852",
          6374 => x"953d7052",
          6375 => x"58d1833f",
          6376 => x"8285ec08",
          6377 => x"558285ec",
          6378 => x"0881dd38",
          6379 => x"0280fb05",
          6380 => x"3370852a",
          6381 => x"70810651",
          6382 => x"55568655",
          6383 => x"7381c938",
          6384 => x"75982b54",
          6385 => x"80742481",
          6386 => x"bf380280",
          6387 => x"d6053370",
          6388 => x"81065854",
          6389 => x"87557681",
          6390 => x"af386b52",
          6391 => x"7851cc9a",
          6392 => x"3f8285ec",
          6393 => x"0874842a",
          6394 => x"70810651",
          6395 => x"55567380",
          6396 => x"2e80d438",
          6397 => x"78548285",
          6398 => x"ec089415",
          6399 => x"082e8188",
          6400 => x"38735a82",
          6401 => x"85ec085c",
          6402 => x"76528a3d",
          6403 => x"705254c7",
          6404 => x"8a3f8285",
          6405 => x"ec085582",
          6406 => x"85ec0880",
          6407 => x"eb388285",
          6408 => x"ec085273",
          6409 => x"51ccba3f",
          6410 => x"8285ec08",
          6411 => x"558285ec",
          6412 => x"08863887",
          6413 => x"5580d139",
          6414 => x"8285ec08",
          6415 => x"842e8838",
          6416 => x"8285ec08",
          6417 => x"80c23877",
          6418 => x"51ce973f",
          6419 => x"8285ec08",
          6420 => x"8285ec08",
          6421 => x"09810570",
          6422 => x"8285ec08",
          6423 => x"07802551",
          6424 => x"55557580",
          6425 => x"2e943873",
          6426 => x"802e8f38",
          6427 => x"80537552",
          6428 => x"7751c0e0",
          6429 => x"3f8285ec",
          6430 => x"0855748c",
          6431 => x"387851ff",
          6432 => x"bac23f82",
          6433 => x"85ec0855",
          6434 => x"748285ec",
          6435 => x"0ca03d0d",
          6436 => x"04e93d0d",
          6437 => x"8253993d",
          6438 => x"c005529a",
          6439 => x"3d51d8b6",
          6440 => x"3f8285ec",
          6441 => x"08548285",
          6442 => x"ec0882b0",
          6443 => x"38785e69",
          6444 => x"528e3d70",
          6445 => x"5258ceea",
          6446 => x"3f8285ec",
          6447 => x"08548285",
          6448 => x"ec088638",
          6449 => x"88548294",
          6450 => x"398285ec",
          6451 => x"08842e09",
          6452 => x"81068288",
          6453 => x"380280df",
          6454 => x"05337085",
          6455 => x"2a810651",
          6456 => x"55865474",
          6457 => x"81f63878",
          6458 => x"5a74528a",
          6459 => x"3d705257",
          6460 => x"c18e3f82",
          6461 => x"85ec0875",
          6462 => x"55568285",
          6463 => x"ec088338",
          6464 => x"87548285",
          6465 => x"ec08812e",
          6466 => x"09810683",
          6467 => x"38825482",
          6468 => x"85ec08ff",
          6469 => x"2e098106",
          6470 => x"86388154",
          6471 => x"81b43973",
          6472 => x"81b03882",
          6473 => x"85ec0852",
          6474 => x"7851c3f5",
          6475 => x"3f8285ec",
          6476 => x"08548285",
          6477 => x"ec08819a",
          6478 => x"388b53a0",
          6479 => x"52b41951",
          6480 => x"ffb6d03f",
          6481 => x"7854ae0b",
          6482 => x"b4153478",
          6483 => x"54900bbf",
          6484 => x"15348288",
          6485 => x"b20a5280",
          6486 => x"ca1951ff",
          6487 => x"b5e33f75",
          6488 => x"5378b411",
          6489 => x"5351c9cb",
          6490 => x"3fa05378",
          6491 => x"b4115380",
          6492 => x"d40551ff",
          6493 => x"b5fa3f78",
          6494 => x"54ae0b80",
          6495 => x"d515347f",
          6496 => x"537880d4",
          6497 => x"115351c9",
          6498 => x"aa3f7854",
          6499 => x"810b8315",
          6500 => x"347751ca",
          6501 => x"f73f8285",
          6502 => x"ec085482",
          6503 => x"85ec08b2",
          6504 => x"388288b2",
          6505 => x"0a526496",
          6506 => x"0551ffb5",
          6507 => x"943f7553",
          6508 => x"64527851",
          6509 => x"c8fd3f64",
          6510 => x"54900b8b",
          6511 => x"15347854",
          6512 => x"810b8315",
          6513 => x"347851ff",
          6514 => x"b7fa3f82",
          6515 => x"85ec0854",
          6516 => x"8b398053",
          6517 => x"75527651",
          6518 => x"ffbdf93f",
          6519 => x"738285ec",
          6520 => x"0c993d0d",
          6521 => x"04da3d0d",
          6522 => x"a93d8405",
          6523 => x"51d2d43f",
          6524 => x"8253a83d",
          6525 => x"ff840552",
          6526 => x"a93d51d5",
          6527 => x"d93f8285",
          6528 => x"ec085582",
          6529 => x"85ec0882",
          6530 => x"d338784d",
          6531 => x"a93d0852",
          6532 => x"9d3d7052",
          6533 => x"58cc8b3f",
          6534 => x"8285ec08",
          6535 => x"558285ec",
          6536 => x"0882b938",
          6537 => x"02819b05",
          6538 => x"3381a006",
          6539 => x"54865573",
          6540 => x"82aa38a0",
          6541 => x"53a43d08",
          6542 => x"52a83dff",
          6543 => x"880551ff",
          6544 => x"b4ae3fac",
          6545 => x"53775292",
          6546 => x"3d705254",
          6547 => x"ffb4a13f",
          6548 => x"aa3d0852",
          6549 => x"7351cbca",
          6550 => x"3f8285ec",
          6551 => x"08558285",
          6552 => x"ec089538",
          6553 => x"636f2e09",
          6554 => x"81068838",
          6555 => x"65a23d08",
          6556 => x"2e923888",
          6557 => x"5581e539",
          6558 => x"8285ec08",
          6559 => x"842e0981",
          6560 => x"0681b838",
          6561 => x"7351c984",
          6562 => x"3f8285ec",
          6563 => x"08558285",
          6564 => x"ec0881c8",
          6565 => x"38685693",
          6566 => x"53a83dff",
          6567 => x"9505528d",
          6568 => x"1651ffb3",
          6569 => x"cb3f02af",
          6570 => x"05338b17",
          6571 => x"348b1633",
          6572 => x"70842a70",
          6573 => x"81065155",
          6574 => x"55738938",
          6575 => x"74a00754",
          6576 => x"738b1734",
          6577 => x"7854810b",
          6578 => x"8315348b",
          6579 => x"16337084",
          6580 => x"2a708106",
          6581 => x"51555573",
          6582 => x"802e80e5",
          6583 => x"386e642e",
          6584 => x"80df3875",
          6585 => x"527851c6",
          6586 => x"913f8285",
          6587 => x"ec085278",
          6588 => x"51ffb6ff",
          6589 => x"3f825582",
          6590 => x"85ec0880",
          6591 => x"2e80dd38",
          6592 => x"8285ec08",
          6593 => x"527851ff",
          6594 => x"b4f33f82",
          6595 => x"85ec0879",
          6596 => x"80d41158",
          6597 => x"58558285",
          6598 => x"ec0880c0",
          6599 => x"38811633",
          6600 => x"5473ae2e",
          6601 => x"09810699",
          6602 => x"38635375",
          6603 => x"527651c6",
          6604 => x"823f7854",
          6605 => x"810b8315",
          6606 => x"34873982",
          6607 => x"85ec089c",
          6608 => x"387751c8",
          6609 => x"9d3f8285",
          6610 => x"ec085582",
          6611 => x"85ec088c",
          6612 => x"387851ff",
          6613 => x"b4ee3f82",
          6614 => x"85ec0855",
          6615 => x"748285ec",
          6616 => x"0ca83d0d",
          6617 => x"04ed3d0d",
          6618 => x"0280db05",
          6619 => x"33028405",
          6620 => x"80df0533",
          6621 => x"57578253",
          6622 => x"953dd005",
          6623 => x"52963d51",
          6624 => x"d2d43f82",
          6625 => x"85ec0855",
          6626 => x"8285ec08",
          6627 => x"80cf3878",
          6628 => x"5a655295",
          6629 => x"3dd40551",
          6630 => x"c9883f82",
          6631 => x"85ec0855",
          6632 => x"8285ec08",
          6633 => x"b8380280",
          6634 => x"cf053381",
          6635 => x"a0065486",
          6636 => x"5573aa38",
          6637 => x"75a70661",
          6638 => x"71098b12",
          6639 => x"3371067a",
          6640 => x"74060751",
          6641 => x"57555674",
          6642 => x"8b153478",
          6643 => x"54810b83",
          6644 => x"15347851",
          6645 => x"ffb3ed3f",
          6646 => x"8285ec08",
          6647 => x"55748285",
          6648 => x"ec0c953d",
          6649 => x"0d04ef3d",
          6650 => x"0d645682",
          6651 => x"53933dd0",
          6652 => x"0552943d",
          6653 => x"51d1df3f",
          6654 => x"8285ec08",
          6655 => x"558285ec",
          6656 => x"0880cb38",
          6657 => x"76586352",
          6658 => x"933dd405",
          6659 => x"51c8933f",
          6660 => x"8285ec08",
          6661 => x"558285ec",
          6662 => x"08b43802",
          6663 => x"80c70533",
          6664 => x"81a00654",
          6665 => x"865573a6",
          6666 => x"38841622",
          6667 => x"86172271",
          6668 => x"902b0753",
          6669 => x"54961f51",
          6670 => x"ffb0863f",
          6671 => x"7654810b",
          6672 => x"83153476",
          6673 => x"51ffb2fc",
          6674 => x"3f8285ec",
          6675 => x"08557482",
          6676 => x"85ec0c93",
          6677 => x"3d0d04ea",
          6678 => x"3d0d696b",
          6679 => x"5c5a8053",
          6680 => x"983dd005",
          6681 => x"52993d51",
          6682 => x"d0ec3f82",
          6683 => x"85ec0882",
          6684 => x"85ec0809",
          6685 => x"81057082",
          6686 => x"85ec0807",
          6687 => x"80255155",
          6688 => x"5779802e",
          6689 => x"81853881",
          6690 => x"70750655",
          6691 => x"5573802e",
          6692 => x"80f9387b",
          6693 => x"5d805f80",
          6694 => x"528d3d70",
          6695 => x"5254ffbd",
          6696 => x"fa3f8285",
          6697 => x"ec085782",
          6698 => x"85ec0880",
          6699 => x"d1387452",
          6700 => x"7351c3ad",
          6701 => x"3f8285ec",
          6702 => x"08578285",
          6703 => x"ec08bf38",
          6704 => x"8285ec08",
          6705 => x"8285ec08",
          6706 => x"655b5956",
          6707 => x"78188119",
          6708 => x"7b185659",
          6709 => x"55743374",
          6710 => x"34811656",
          6711 => x"8a7827ec",
          6712 => x"388b5675",
          6713 => x"1a548074",
          6714 => x"3475802e",
          6715 => x"9e38ff16",
          6716 => x"701b7033",
          6717 => x"51555673",
          6718 => x"a02ee838",
          6719 => x"8e397684",
          6720 => x"2e098106",
          6721 => x"8638807a",
          6722 => x"34805776",
          6723 => x"09810570",
          6724 => x"78078025",
          6725 => x"51547a80",
          6726 => x"2e80c138",
          6727 => x"73802ebc",
          6728 => x"387ba011",
          6729 => x"085351ff",
          6730 => x"b0d33f82",
          6731 => x"85ec0857",
          6732 => x"8285ec08",
          6733 => x"a7387b70",
          6734 => x"33555580",
          6735 => x"c3567383",
          6736 => x"2e8b3880",
          6737 => x"e4567384",
          6738 => x"2e8338a7",
          6739 => x"567515b4",
          6740 => x"0551ffad",
          6741 => x"a33f8285",
          6742 => x"ec087b0c",
          6743 => x"768285ec",
          6744 => x"0c983d0d",
          6745 => x"04e63d0d",
          6746 => x"82539c3d",
          6747 => x"ffb80552",
          6748 => x"9d3d51ce",
          6749 => x"e13f8285",
          6750 => x"ec088285",
          6751 => x"ec085654",
          6752 => x"8285ec08",
          6753 => x"8398388b",
          6754 => x"53a0528b",
          6755 => x"3d705259",
          6756 => x"ffae803f",
          6757 => x"736d7033",
          6758 => x"7081ff06",
          6759 => x"52575557",
          6760 => x"9f742781",
          6761 => x"bc387858",
          6762 => x"7481ff06",
          6763 => x"6d81054e",
          6764 => x"705255ff",
          6765 => x"aec93f82",
          6766 => x"85ec0880",
          6767 => x"2ea5386c",
          6768 => x"70337053",
          6769 => x"5754ffae",
          6770 => x"bd3f8285",
          6771 => x"ec08802e",
          6772 => x"8d387488",
          6773 => x"2b76076d",
          6774 => x"81054e55",
          6775 => x"86398285",
          6776 => x"ec0855ff",
          6777 => x"9f157083",
          6778 => x"ffff0651",
          6779 => x"54739926",
          6780 => x"8a38e015",
          6781 => x"7083ffff",
          6782 => x"06565480",
          6783 => x"ff752787",
          6784 => x"3881feb4",
          6785 => x"15335574",
          6786 => x"802ea338",
          6787 => x"74528280",
          6788 => x"b451ffad",
          6789 => x"c93f8285",
          6790 => x"ec089338",
          6791 => x"81ff7527",
          6792 => x"88387689",
          6793 => x"2688388b",
          6794 => x"398a7727",
          6795 => x"86388655",
          6796 => x"81ec3981",
          6797 => x"ff75278f",
          6798 => x"3874882a",
          6799 => x"54737870",
          6800 => x"81055a34",
          6801 => x"81175774",
          6802 => x"78708105",
          6803 => x"5a348117",
          6804 => x"6d703370",
          6805 => x"81ff0652",
          6806 => x"57555773",
          6807 => x"9f26fec8",
          6808 => x"388b3d33",
          6809 => x"54865573",
          6810 => x"81e52e81",
          6811 => x"b1387680",
          6812 => x"2e993802",
          6813 => x"a7055576",
          6814 => x"15703351",
          6815 => x"5473a02e",
          6816 => x"09810687",
          6817 => x"38ff1757",
          6818 => x"76ed3879",
          6819 => x"41804380",
          6820 => x"52913d70",
          6821 => x"5255ffba",
          6822 => x"823f8285",
          6823 => x"ec085482",
          6824 => x"85ec0880",
          6825 => x"f7388152",
          6826 => x"7451ffbf",
          6827 => x"b43f8285",
          6828 => x"ec085482",
          6829 => x"85ec088d",
          6830 => x"387680c4",
          6831 => x"386754e5",
          6832 => x"743480c6",
          6833 => x"398285ec",
          6834 => x"08842e09",
          6835 => x"810680cc",
          6836 => x"38805476",
          6837 => x"742e80c4",
          6838 => x"38815274",
          6839 => x"51ffbcff",
          6840 => x"3f8285ec",
          6841 => x"08548285",
          6842 => x"ec08b138",
          6843 => x"a0538285",
          6844 => x"ec085267",
          6845 => x"51ffab9b",
          6846 => x"3f675488",
          6847 => x"0b8b1534",
          6848 => x"8b537852",
          6849 => x"6751ffaa",
          6850 => x"e73f7954",
          6851 => x"810b8315",
          6852 => x"347951ff",
          6853 => x"adae3f82",
          6854 => x"85ec0854",
          6855 => x"73557482",
          6856 => x"85ec0c9c",
          6857 => x"3d0d04f2",
          6858 => x"3d0d6062",
          6859 => x"02880580",
          6860 => x"cb053393",
          6861 => x"3dfc0555",
          6862 => x"7254405e",
          6863 => x"5ad2c83f",
          6864 => x"8285ec08",
          6865 => x"588285ec",
          6866 => x"0882bf38",
          6867 => x"911a3358",
          6868 => x"7782b738",
          6869 => x"7c802e97",
          6870 => x"388c1a08",
          6871 => x"59789038",
          6872 => x"901a3370",
          6873 => x"812a7081",
          6874 => x"06515555",
          6875 => x"73903887",
          6876 => x"54829939",
          6877 => x"82588292",
          6878 => x"39815882",
          6879 => x"8d397e8a",
          6880 => x"11227089",
          6881 => x"2b70557f",
          6882 => x"54565656",
          6883 => x"fec6fb3f",
          6884 => x"ff147d06",
          6885 => x"70098105",
          6886 => x"7072079f",
          6887 => x"2a8285ec",
          6888 => x"08058c19",
          6889 => x"087c405a",
          6890 => x"5d555581",
          6891 => x"77278838",
          6892 => x"98160877",
          6893 => x"26833882",
          6894 => x"57767756",
          6895 => x"59805674",
          6896 => x"527951ff",
          6897 => x"adde3f81",
          6898 => x"157f5555",
          6899 => x"98140875",
          6900 => x"26833882",
          6901 => x"558285ec",
          6902 => x"08812eff",
          6903 => x"97388285",
          6904 => x"ec08ff2e",
          6905 => x"ff933882",
          6906 => x"85ec088e",
          6907 => x"38811656",
          6908 => x"757b2e09",
          6909 => x"81068738",
          6910 => x"93397459",
          6911 => x"80567477",
          6912 => x"2e098106",
          6913 => x"ffb93887",
          6914 => x"5880ff39",
          6915 => x"7d802eba",
          6916 => x"38787b55",
          6917 => x"557a802e",
          6918 => x"b4388115",
          6919 => x"5673812e",
          6920 => x"09810683",
          6921 => x"38ff5675",
          6922 => x"5374527e",
          6923 => x"51ffaeed",
          6924 => x"3f8285ec",
          6925 => x"08588285",
          6926 => x"ec0880ce",
          6927 => x"38748116",
          6928 => x"ff165656",
          6929 => x"5c73d338",
          6930 => x"8439ff19",
          6931 => x"5c7e7c8c",
          6932 => x"120c557d",
          6933 => x"802eb338",
          6934 => x"78881b0c",
          6935 => x"7c8c1b0c",
          6936 => x"901a3380",
          6937 => x"c0075473",
          6938 => x"901b3498",
          6939 => x"1508fe05",
          6940 => x"90160857",
          6941 => x"54757426",
          6942 => x"9138757b",
          6943 => x"3190160c",
          6944 => x"84153381",
          6945 => x"07547384",
          6946 => x"16347754",
          6947 => x"738285ec",
          6948 => x"0c903d0d",
          6949 => x"04e93d0d",
          6950 => x"6b6d0288",
          6951 => x"0580eb05",
          6952 => x"339d3d54",
          6953 => x"5a5c59c5",
          6954 => x"9a3f8b56",
          6955 => x"800b8285",
          6956 => x"ec08248c",
          6957 => x"82388285",
          6958 => x"ec08822b",
          6959 => x"829d9011",
          6960 => x"08515574",
          6961 => x"802e8438",
          6962 => x"80753482",
          6963 => x"85ec0881",
          6964 => x"ff065f81",
          6965 => x"527e51ff",
          6966 => x"a08f3f82",
          6967 => x"85ec0881",
          6968 => x"ff067081",
          6969 => x"06565783",
          6970 => x"56748bcb",
          6971 => x"3876822a",
          6972 => x"70810651",
          6973 => x"558a5674",
          6974 => x"8bbd3899",
          6975 => x"3dfc0553",
          6976 => x"83527e51",
          6977 => x"ffa4af3f",
          6978 => x"8285ec08",
          6979 => x"99386755",
          6980 => x"74802e92",
          6981 => x"38748280",
          6982 => x"80268b38",
          6983 => x"ff157506",
          6984 => x"5574802e",
          6985 => x"83388148",
          6986 => x"78802e87",
          6987 => x"38848079",
          6988 => x"26923878",
          6989 => x"81800a26",
          6990 => x"8b38ff19",
          6991 => x"79065574",
          6992 => x"802e8638",
          6993 => x"93568aef",
          6994 => x"3978892a",
          6995 => x"6e892a70",
          6996 => x"892b7759",
          6997 => x"4843597a",
          6998 => x"83388156",
          6999 => x"61098105",
          7000 => x"70802577",
          7001 => x"07515591",
          7002 => x"56748acb",
          7003 => x"38993df8",
          7004 => x"05538152",
          7005 => x"7e51ffa3",
          7006 => x"bd3f8156",
          7007 => x"8285ec08",
          7008 => x"8ab53877",
          7009 => x"832a7077",
          7010 => x"068285ec",
          7011 => x"08435645",
          7012 => x"748338bf",
          7013 => x"4166558e",
          7014 => x"56607526",
          7015 => x"8a993874",
          7016 => x"61317048",
          7017 => x"5580ff75",
          7018 => x"278a8c38",
          7019 => x"93567881",
          7020 => x"80268a83",
          7021 => x"3877812a",
          7022 => x"70810656",
          7023 => x"4374802e",
          7024 => x"95387787",
          7025 => x"06557482",
          7026 => x"2e839438",
          7027 => x"77810655",
          7028 => x"74802e83",
          7029 => x"8a387781",
          7030 => x"06559356",
          7031 => x"825e7480",
          7032 => x"2e89d438",
          7033 => x"785a7d83",
          7034 => x"2e098106",
          7035 => x"80e03878",
          7036 => x"ae386691",
          7037 => x"2a57810b",
          7038 => x"8280d822",
          7039 => x"565a7480",
          7040 => x"2e9d3874",
          7041 => x"77269838",
          7042 => x"8280d856",
          7043 => x"79108217",
          7044 => x"70225757",
          7045 => x"5a74802e",
          7046 => x"86387675",
          7047 => x"27ee3879",
          7048 => x"526651fe",
          7049 => x"c1e43f82",
          7050 => x"85ec0882",
          7051 => x"2b848711",
          7052 => x"892a5e55",
          7053 => x"a05c800b",
          7054 => x"8285ec08",
          7055 => x"fc808a05",
          7056 => x"5644fdff",
          7057 => x"f00a7527",
          7058 => x"80f23888",
          7059 => x"dd3978ae",
          7060 => x"38668c2a",
          7061 => x"57810b82",
          7062 => x"80c82256",
          7063 => x"5a74802e",
          7064 => x"9d387477",
          7065 => x"26983882",
          7066 => x"80c85679",
          7067 => x"10821770",
          7068 => x"2257575a",
          7069 => x"74802e86",
          7070 => x"38767527",
          7071 => x"ee387952",
          7072 => x"6651fec1",
          7073 => x"853f8285",
          7074 => x"ec088285",
          7075 => x"ec080584",
          7076 => x"05578285",
          7077 => x"ec089ff5",
          7078 => x"26983881",
          7079 => x"0b8285ec",
          7080 => x"08712b82",
          7081 => x"85ec0811",
          7082 => x"1270732a",
          7083 => x"83055a51",
          7084 => x"565e83ff",
          7085 => x"17892a5d",
          7086 => x"815ca044",
          7087 => x"601c7d11",
          7088 => x"65056970",
          7089 => x"12ff0571",
          7090 => x"09810570",
          7091 => x"72067431",
          7092 => x"5c525957",
          7093 => x"59407d83",
          7094 => x"2e098106",
          7095 => x"8938761c",
          7096 => x"6018415c",
          7097 => x"8439761d",
          7098 => x"5d79842b",
          7099 => x"70196231",
          7100 => x"68585155",
          7101 => x"74762687",
          7102 => x"b138757c",
          7103 => x"317d317a",
          7104 => x"53706531",
          7105 => x"5255fec0",
          7106 => x"813f8285",
          7107 => x"ec08587d",
          7108 => x"832e0981",
          7109 => x"069b3882",
          7110 => x"85ec0883",
          7111 => x"fff52680",
          7112 => x"dd387887",
          7113 => x"85387981",
          7114 => x"2a5978fd",
          7115 => x"b73886fa",
          7116 => x"397d822e",
          7117 => x"09810680",
          7118 => x"c53883ff",
          7119 => x"f50b8285",
          7120 => x"ec0827a0",
          7121 => x"38788f38",
          7122 => x"791a5574",
          7123 => x"80c02686",
          7124 => x"387459fd",
          7125 => x"8f396281",
          7126 => x"06557480",
          7127 => x"2e8f3883",
          7128 => x"5efd8139",
          7129 => x"8285ec08",
          7130 => x"9ff52692",
          7131 => x"387886ba",
          7132 => x"38791a59",
          7133 => x"81807927",
          7134 => x"fcea3886",
          7135 => x"ad398055",
          7136 => x"7d812e09",
          7137 => x"81068338",
          7138 => x"7d559ff5",
          7139 => x"78278b38",
          7140 => x"74810655",
          7141 => x"8e567486",
          7142 => x"9e388480",
          7143 => x"5380527a",
          7144 => x"51ffa1ef",
          7145 => x"3f8b5381",
          7146 => x"fef0527a",
          7147 => x"51ffa1c0",
          7148 => x"3f848052",
          7149 => x"8b1b51ff",
          7150 => x"a0e93f79",
          7151 => x"8d1c347b",
          7152 => x"83ffff06",
          7153 => x"528e1b51",
          7154 => x"ffa0d83f",
          7155 => x"810b901c",
          7156 => x"347d8332",
          7157 => x"70098105",
          7158 => x"70962a84",
          7159 => x"80065451",
          7160 => x"55911b51",
          7161 => x"ffa0bc3f",
          7162 => x"66557483",
          7163 => x"ffff2690",
          7164 => x"387483ff",
          7165 => x"ff065293",
          7166 => x"1b51ffa0",
          7167 => x"a63f8a39",
          7168 => x"7452a01b",
          7169 => x"51ffa0b9",
          7170 => x"3ff80b95",
          7171 => x"1c34bf52",
          7172 => x"981b51ff",
          7173 => x"a08d3f81",
          7174 => x"ff529a1b",
          7175 => x"51ffa083",
          7176 => x"3f60529c",
          7177 => x"1b51ffa0",
          7178 => x"983f7d83",
          7179 => x"2e098106",
          7180 => x"80cb3882",
          7181 => x"88b20a52",
          7182 => x"80c31b51",
          7183 => x"ffa0823f",
          7184 => x"7c52a41b",
          7185 => x"51ff9ff9",
          7186 => x"3f8252ac",
          7187 => x"1b51ff9f",
          7188 => x"f03f8152",
          7189 => x"b01b51ff",
          7190 => x"9fc93f86",
          7191 => x"52b21b51",
          7192 => x"ff9fc03f",
          7193 => x"ff800b80",
          7194 => x"c01c34a9",
          7195 => x"0b80c21c",
          7196 => x"34935381",
          7197 => x"fefc5280",
          7198 => x"c71b51ae",
          7199 => x"398288b2",
          7200 => x"0a52a71b",
          7201 => x"51ff9fb9",
          7202 => x"3f7c83ff",
          7203 => x"ff065296",
          7204 => x"1b51ff9f",
          7205 => x"8e3fff80",
          7206 => x"0ba41c34",
          7207 => x"a90ba61c",
          7208 => x"34935381",
          7209 => x"ff9052ab",
          7210 => x"1b51ff9f",
          7211 => x"c33f82d4",
          7212 => x"d55283fe",
          7213 => x"1b705259",
          7214 => x"ff9ee83f",
          7215 => x"81546053",
          7216 => x"7a527e51",
          7217 => x"ff9b8b3f",
          7218 => x"81568285",
          7219 => x"ec0883e7",
          7220 => x"387d832e",
          7221 => x"09810680",
          7222 => x"ee387554",
          7223 => x"60860553",
          7224 => x"7a527e51",
          7225 => x"ff9aeb3f",
          7226 => x"84805380",
          7227 => x"527a51ff",
          7228 => x"9fa13f84",
          7229 => x"8b85a4d2",
          7230 => x"527a51ff",
          7231 => x"9ec33f86",
          7232 => x"8a85e4f2",
          7233 => x"5283e41b",
          7234 => x"51ff9eb5",
          7235 => x"3fff1852",
          7236 => x"83e81b51",
          7237 => x"ff9eaa3f",
          7238 => x"825283ec",
          7239 => x"1b51ff9e",
          7240 => x"a03f82d4",
          7241 => x"d5527851",
          7242 => x"ff9df83f",
          7243 => x"75546087",
          7244 => x"05537a52",
          7245 => x"7e51ff9a",
          7246 => x"993f7554",
          7247 => x"6016537a",
          7248 => x"527e51ff",
          7249 => x"9a8c3f65",
          7250 => x"5380527a",
          7251 => x"51ff9ec3",
          7252 => x"3f7f5680",
          7253 => x"587d832e",
          7254 => x"0981069a",
          7255 => x"38f8527a",
          7256 => x"51ff9ddd",
          7257 => x"3fff5284",
          7258 => x"1b51ff9d",
          7259 => x"d43ff00a",
          7260 => x"52881b51",
          7261 => x"913987ff",
          7262 => x"fff8557d",
          7263 => x"812e8338",
          7264 => x"f8557452",
          7265 => x"7a51ff9d",
          7266 => x"b83f7c55",
          7267 => x"61577462",
          7268 => x"26833874",
          7269 => x"57765475",
          7270 => x"537a527e",
          7271 => x"51ff99b2",
          7272 => x"3f8285ec",
          7273 => x"08828738",
          7274 => x"84805382",
          7275 => x"85ec0852",
          7276 => x"7a51ff9d",
          7277 => x"de3f7616",
          7278 => x"75783156",
          7279 => x"5674cd38",
          7280 => x"81185877",
          7281 => x"802eff8d",
          7282 => x"3879557d",
          7283 => x"832e8338",
          7284 => x"63556157",
          7285 => x"74622683",
          7286 => x"38745776",
          7287 => x"5475537a",
          7288 => x"527e51ff",
          7289 => x"98ec3f82",
          7290 => x"85ec0881",
          7291 => x"c1387616",
          7292 => x"75783156",
          7293 => x"5674db38",
          7294 => x"8c567d83",
          7295 => x"2e933886",
          7296 => x"566683ff",
          7297 => x"ff268a38",
          7298 => x"84567d82",
          7299 => x"2e833881",
          7300 => x"56648106",
          7301 => x"587780fe",
          7302 => x"38848053",
          7303 => x"77527a51",
          7304 => x"ff9cf03f",
          7305 => x"82d4d552",
          7306 => x"7851ff9b",
          7307 => x"f63f83be",
          7308 => x"1b557775",
          7309 => x"34810b81",
          7310 => x"1634810b",
          7311 => x"82163477",
          7312 => x"83163475",
          7313 => x"84163460",
          7314 => x"67055680",
          7315 => x"fdc15275",
          7316 => x"51feb9b6",
          7317 => x"3ffe0b85",
          7318 => x"16348285",
          7319 => x"ec08822a",
          7320 => x"bf075675",
          7321 => x"86163482",
          7322 => x"85ec0887",
          7323 => x"16346052",
          7324 => x"83c61b51",
          7325 => x"ff9bca3f",
          7326 => x"665283ca",
          7327 => x"1b51ff9b",
          7328 => x"c03f8154",
          7329 => x"77537a52",
          7330 => x"7e51ff97",
          7331 => x"c53f8156",
          7332 => x"8285ec08",
          7333 => x"a2388053",
          7334 => x"80527e51",
          7335 => x"ff99973f",
          7336 => x"81568285",
          7337 => x"ec089038",
          7338 => x"89398e56",
          7339 => x"8a398156",
          7340 => x"86398285",
          7341 => x"ec085675",
          7342 => x"8285ec0c",
          7343 => x"993d0d04",
          7344 => x"f53d0d7d",
          7345 => x"605b5980",
          7346 => x"7960ff05",
          7347 => x"5a575776",
          7348 => x"7825b438",
          7349 => x"8d3df811",
          7350 => x"55558153",
          7351 => x"fc155279",
          7352 => x"51c9c03f",
          7353 => x"7a812e09",
          7354 => x"81069c38",
          7355 => x"8c3d3355",
          7356 => x"748d2edb",
          7357 => x"38747670",
          7358 => x"81055834",
          7359 => x"81175774",
          7360 => x"8a2e0981",
          7361 => x"06c93880",
          7362 => x"76347855",
          7363 => x"76833876",
          7364 => x"55748285",
          7365 => x"ec0c8d3d",
          7366 => x"0d04f73d",
          7367 => x"0d7b0284",
          7368 => x"05b30533",
          7369 => x"5957778a",
          7370 => x"2e098106",
          7371 => x"87388d52",
          7372 => x"7651e73f",
          7373 => x"84170856",
          7374 => x"80762480",
          7375 => x"c2388817",
          7376 => x"0877178c",
          7377 => x"05565977",
          7378 => x"75348116",
          7379 => x"56bb7625",
          7380 => x"a5388b3d",
          7381 => x"fc055475",
          7382 => x"538c1752",
          7383 => x"760851cb",
          7384 => x"bf3f7976",
          7385 => x"32700981",
          7386 => x"05707207",
          7387 => x"9f2a7009",
          7388 => x"81055351",
          7389 => x"56567584",
          7390 => x"180c8119",
          7391 => x"88180c8b",
          7392 => x"3d0d04f9",
          7393 => x"3d0d7984",
          7394 => x"11085656",
          7395 => x"807524a7",
          7396 => x"38893dfc",
          7397 => x"05547453",
          7398 => x"8c165275",
          7399 => x"0851cb80",
          7400 => x"3f8285ec",
          7401 => x"08913884",
          7402 => x"1608782e",
          7403 => x"09810687",
          7404 => x"38881608",
          7405 => x"558339ff",
          7406 => x"55748285",
          7407 => x"ec0c893d",
          7408 => x"0d04fd3d",
          7409 => x"0d755480",
          7410 => x"cc538052",
          7411 => x"7351ff99",
          7412 => x"c23f7674",
          7413 => x"0c853d0d",
          7414 => x"04ea3d0d",
          7415 => x"0280e305",
          7416 => x"336a5386",
          7417 => x"3d705354",
          7418 => x"54d83f73",
          7419 => x"527251fe",
          7420 => x"a93f7251",
          7421 => x"ff8d3f98",
          7422 => x"3d0d0400",
          7423 => x"00ffffff",
          7424 => x"ff00ffff",
          7425 => x"ffff00ff",
          7426 => x"ffffff00",
          7427 => x"0000118e",
          7428 => x"00001112",
          7429 => x"00001119",
          7430 => x"00001120",
          7431 => x"00001127",
          7432 => x"0000112e",
          7433 => x"00001135",
          7434 => x"0000113c",
          7435 => x"00001143",
          7436 => x"0000114a",
          7437 => x"00001151",
          7438 => x"00001158",
          7439 => x"0000115e",
          7440 => x"00001164",
          7441 => x"0000116a",
          7442 => x"00001170",
          7443 => x"00001176",
          7444 => x"0000117c",
          7445 => x"00001182",
          7446 => x"00001188",
          7447 => x"000026ce",
          7448 => x"000026d4",
          7449 => x"000026da",
          7450 => x"000026e0",
          7451 => x"000026e6",
          7452 => x"000032e6",
          7453 => x"000033d0",
          7454 => x"000034bd",
          7455 => x"000036eb",
          7456 => x"000033b8",
          7457 => x"000031c3",
          7458 => x"00003567",
          7459 => x"000036c2",
          7460 => x"000035a4",
          7461 => x"0000363b",
          7462 => x"000035c0",
          7463 => x"0000346d",
          7464 => x"000031c3",
          7465 => x"000034bd",
          7466 => x"000034e0",
          7467 => x"00003567",
          7468 => x"000031c3",
          7469 => x"000031c3",
          7470 => x"000035c0",
          7471 => x"0000363b",
          7472 => x"000036c2",
          7473 => x"000036eb",
          7474 => x"64696e69",
          7475 => x"74000000",
          7476 => x"64696f63",
          7477 => x"746c0000",
          7478 => x"66696e69",
          7479 => x"74000000",
          7480 => x"666c6f61",
          7481 => x"64000000",
          7482 => x"66657865",
          7483 => x"63000000",
          7484 => x"6d636c65",
          7485 => x"61720000",
          7486 => x"6d636f70",
          7487 => x"79000000",
          7488 => x"6d646966",
          7489 => x"66000000",
          7490 => x"6d64756d",
          7491 => x"70000000",
          7492 => x"6d656200",
          7493 => x"6d656800",
          7494 => x"6d657700",
          7495 => x"68696400",
          7496 => x"68696500",
          7497 => x"68666400",
          7498 => x"68666500",
          7499 => x"63616c6c",
          7500 => x"00000000",
          7501 => x"6a6d7000",
          7502 => x"72657374",
          7503 => x"61727400",
          7504 => x"72657365",
          7505 => x"74000000",
          7506 => x"696e666f",
          7507 => x"00000000",
          7508 => x"74657374",
          7509 => x"00000000",
          7510 => x"74626173",
          7511 => x"69630000",
          7512 => x"6d626173",
          7513 => x"69630000",
          7514 => x"6b696c6f",
          7515 => x"00000000",
          7516 => x"65640000",
          7517 => x"4469736b",
          7518 => x"20457272",
          7519 => x"6f720a00",
          7520 => x"496e7465",
          7521 => x"726e616c",
          7522 => x"20657272",
          7523 => x"6f722e0a",
          7524 => x"00000000",
          7525 => x"4469736b",
          7526 => x"206e6f74",
          7527 => x"20726561",
          7528 => x"64792e0a",
          7529 => x"00000000",
          7530 => x"4e6f2066",
          7531 => x"696c6520",
          7532 => x"666f756e",
          7533 => x"642e0a00",
          7534 => x"4e6f2070",
          7535 => x"61746820",
          7536 => x"666f756e",
          7537 => x"642e0a00",
          7538 => x"496e7661",
          7539 => x"6c696420",
          7540 => x"66696c65",
          7541 => x"6e616d65",
          7542 => x"2e0a0000",
          7543 => x"41636365",
          7544 => x"73732064",
          7545 => x"656e6965",
          7546 => x"642e0a00",
          7547 => x"46696c65",
          7548 => x"20616c72",
          7549 => x"65616479",
          7550 => x"20657869",
          7551 => x"7374732e",
          7552 => x"0a000000",
          7553 => x"46696c65",
          7554 => x"2068616e",
          7555 => x"646c6520",
          7556 => x"696e7661",
          7557 => x"6c69642e",
          7558 => x"0a000000",
          7559 => x"53442069",
          7560 => x"73207772",
          7561 => x"69746520",
          7562 => x"70726f74",
          7563 => x"65637465",
          7564 => x"642e0a00",
          7565 => x"44726976",
          7566 => x"65206e75",
          7567 => x"6d626572",
          7568 => x"20697320",
          7569 => x"696e7661",
          7570 => x"6c69642e",
          7571 => x"0a000000",
          7572 => x"4469736b",
          7573 => x"206e6f74",
          7574 => x"20656e61",
          7575 => x"626c6564",
          7576 => x"2e0a0000",
          7577 => x"4e6f2063",
          7578 => x"6f6d7061",
          7579 => x"7469626c",
          7580 => x"65206669",
          7581 => x"6c657379",
          7582 => x"7374656d",
          7583 => x"20666f75",
          7584 => x"6e64206f",
          7585 => x"6e206469",
          7586 => x"736b2e0a",
          7587 => x"00000000",
          7588 => x"466f726d",
          7589 => x"61742061",
          7590 => x"626f7274",
          7591 => x"65642e0a",
          7592 => x"00000000",
          7593 => x"54696d65",
          7594 => x"6f75742c",
          7595 => x"206f7065",
          7596 => x"72617469",
          7597 => x"6f6e2063",
          7598 => x"616e6365",
          7599 => x"6c6c6564",
          7600 => x"2e0a0000",
          7601 => x"46696c65",
          7602 => x"20697320",
          7603 => x"6c6f636b",
          7604 => x"65642e0a",
          7605 => x"00000000",
          7606 => x"496e7375",
          7607 => x"66666963",
          7608 => x"69656e74",
          7609 => x"206d656d",
          7610 => x"6f72792e",
          7611 => x"0a000000",
          7612 => x"546f6f20",
          7613 => x"6d616e79",
          7614 => x"206f7065",
          7615 => x"6e206669",
          7616 => x"6c65732e",
          7617 => x"0a000000",
          7618 => x"50617261",
          7619 => x"6d657465",
          7620 => x"72732069",
          7621 => x"6e636f72",
          7622 => x"72656374",
          7623 => x"2e0a0000",
          7624 => x"53756363",
          7625 => x"6573732e",
          7626 => x"0a000000",
          7627 => x"556e6b6e",
          7628 => x"6f776e20",
          7629 => x"6572726f",
          7630 => x"722e0a00",
          7631 => x"0a256c75",
          7632 => x"20627974",
          7633 => x"65732025",
          7634 => x"73206174",
          7635 => x"20256c75",
          7636 => x"20627974",
          7637 => x"65732f73",
          7638 => x"65632e0a",
          7639 => x"00000000",
          7640 => x"72656164",
          7641 => x"00000000",
          7642 => x"25303858",
          7643 => x"00000000",
          7644 => x"3a202000",
          7645 => x"25303458",
          7646 => x"00000000",
          7647 => x"20202020",
          7648 => x"20202020",
          7649 => x"00000000",
          7650 => x"25303258",
          7651 => x"00000000",
          7652 => x"20200000",
          7653 => x"207c0000",
          7654 => x"7c0d0a00",
          7655 => x"7a4f5300",
          7656 => x"0a2a2a20",
          7657 => x"25732028",
          7658 => x"00000000",
          7659 => x"30322f30",
          7660 => x"352f3230",
          7661 => x"32300000",
          7662 => x"76312e30",
          7663 => x"32000000",
          7664 => x"205a5055",
          7665 => x"2c207265",
          7666 => x"76202530",
          7667 => x"32782920",
          7668 => x"25732025",
          7669 => x"73202a2a",
          7670 => x"0a0a0000",
          7671 => x"5a505520",
          7672 => x"496e7465",
          7673 => x"72727570",
          7674 => x"74204861",
          7675 => x"6e646c65",
          7676 => x"720a0000",
          7677 => x"54696d65",
          7678 => x"7220696e",
          7679 => x"74657272",
          7680 => x"7570740a",
          7681 => x"00000000",
          7682 => x"50533220",
          7683 => x"696e7465",
          7684 => x"72727570",
          7685 => x"740a0000",
          7686 => x"494f4354",
          7687 => x"4c205244",
          7688 => x"20696e74",
          7689 => x"65727275",
          7690 => x"70740a00",
          7691 => x"494f4354",
          7692 => x"4c205752",
          7693 => x"20696e74",
          7694 => x"65727275",
          7695 => x"70740a00",
          7696 => x"55415254",
          7697 => x"30205258",
          7698 => x"20696e74",
          7699 => x"65727275",
          7700 => x"70740a00",
          7701 => x"55415254",
          7702 => x"30205458",
          7703 => x"20696e74",
          7704 => x"65727275",
          7705 => x"70740a00",
          7706 => x"55415254",
          7707 => x"31205258",
          7708 => x"20696e74",
          7709 => x"65727275",
          7710 => x"70740a00",
          7711 => x"55415254",
          7712 => x"31205458",
          7713 => x"20696e74",
          7714 => x"65727275",
          7715 => x"70740a00",
          7716 => x"53657474",
          7717 => x"696e6720",
          7718 => x"75702074",
          7719 => x"696d6572",
          7720 => x"2e2e2e0a",
          7721 => x"00000000",
          7722 => x"456e6162",
          7723 => x"6c696e67",
          7724 => x"2074696d",
          7725 => x"65722e2e",
          7726 => x"2e0a0000",
          7727 => x"6175746f",
          7728 => x"65786563",
          7729 => x"2e626174",
          7730 => x"00000000",
          7731 => x"7a4f532e",
          7732 => x"68737400",
          7733 => x"303a0000",
          7734 => x"4661696c",
          7735 => x"65642074",
          7736 => x"6f20696e",
          7737 => x"69746961",
          7738 => x"6c697365",
          7739 => x"20736420",
          7740 => x"63617264",
          7741 => x"20302c20",
          7742 => x"706c6561",
          7743 => x"73652069",
          7744 => x"6e697420",
          7745 => x"6d616e75",
          7746 => x"616c6c79",
          7747 => x"2e0a0000",
          7748 => x"2a200000",
          7749 => x"436c6561",
          7750 => x"72696e67",
          7751 => x"2e2e2e2e",
          7752 => x"00000000",
          7753 => x"436f7079",
          7754 => x"696e672e",
          7755 => x"2e2e0000",
          7756 => x"436f6d70",
          7757 => x"6172696e",
          7758 => x"672e2e2e",
          7759 => x"00000000",
          7760 => x"2530386c",
          7761 => x"78282530",
          7762 => x"3878292d",
          7763 => x"3e253038",
          7764 => x"6c782825",
          7765 => x"30387829",
          7766 => x"0a000000",
          7767 => x"44756d70",
          7768 => x"204d656d",
          7769 => x"6f72790a",
          7770 => x"00000000",
          7771 => x"0a436f6d",
          7772 => x"706c6574",
          7773 => x"652e0a00",
          7774 => x"25303858",
          7775 => x"20253032",
          7776 => x"582d0000",
          7777 => x"3f3f3f0a",
          7778 => x"00000000",
          7779 => x"25303858",
          7780 => x"20253034",
          7781 => x"582d0000",
          7782 => x"25303858",
          7783 => x"20253038",
          7784 => x"582d0000",
          7785 => x"45786563",
          7786 => x"7574696e",
          7787 => x"6720636f",
          7788 => x"64652040",
          7789 => x"20253038",
          7790 => x"78202e2e",
          7791 => x"2e0a0000",
          7792 => x"43616c6c",
          7793 => x"696e6720",
          7794 => x"636f6465",
          7795 => x"20402025",
          7796 => x"30387820",
          7797 => x"2e2e2e0a",
          7798 => x"00000000",
          7799 => x"43616c6c",
          7800 => x"20726574",
          7801 => x"75726e65",
          7802 => x"6420636f",
          7803 => x"64652028",
          7804 => x"2564292e",
          7805 => x"0a000000",
          7806 => x"52657374",
          7807 => x"61727469",
          7808 => x"6e672061",
          7809 => x"70706c69",
          7810 => x"63617469",
          7811 => x"6f6e2e2e",
          7812 => x"2e0a0000",
          7813 => x"436f6c64",
          7814 => x"20726562",
          7815 => x"6f6f7469",
          7816 => x"6e672e2e",
          7817 => x"2e0a0000",
          7818 => x"5a505500",
          7819 => x"62696e00",
          7820 => x"25643a5c",
          7821 => x"25735c25",
          7822 => x"732e2573",
          7823 => x"00000000",
          7824 => x"25643a5c",
          7825 => x"25735c25",
          7826 => x"73000000",
          7827 => x"25643a5c",
          7828 => x"25730000",
          7829 => x"42616420",
          7830 => x"636f6d6d",
          7831 => x"616e642e",
          7832 => x"0a000000",
          7833 => x"52756e6e",
          7834 => x"696e672e",
          7835 => x"2e2e0a00",
          7836 => x"456e6162",
          7837 => x"6c696e67",
          7838 => x"20696e74",
          7839 => x"65727275",
          7840 => x"7074732e",
          7841 => x"2e2e0a00",
          7842 => x"25642f25",
          7843 => x"642f2564",
          7844 => x"2025643a",
          7845 => x"25643a25",
          7846 => x"642e2564",
          7847 => x"25640a00",
          7848 => x"536f4320",
          7849 => x"436f6e66",
          7850 => x"69677572",
          7851 => x"6174696f",
          7852 => x"6e000000",
          7853 => x"20286672",
          7854 => x"6f6d2053",
          7855 => x"6f432063",
          7856 => x"6f6e6669",
          7857 => x"67290000",
          7858 => x"3a0a4465",
          7859 => x"76696365",
          7860 => x"7320696d",
          7861 => x"706c656d",
          7862 => x"656e7465",
          7863 => x"643a0a00",
          7864 => x"20202020",
          7865 => x"57422053",
          7866 => x"4452414d",
          7867 => x"20202825",
          7868 => x"3038583a",
          7869 => x"25303858",
          7870 => x"292e0a00",
          7871 => x"20202020",
          7872 => x"53445241",
          7873 => x"4d202020",
          7874 => x"20202825",
          7875 => x"3038583a",
          7876 => x"25303858",
          7877 => x"292e0a00",
          7878 => x"20202020",
          7879 => x"494e534e",
          7880 => x"20425241",
          7881 => x"4d202825",
          7882 => x"3038583a",
          7883 => x"25303858",
          7884 => x"292e0a00",
          7885 => x"20202020",
          7886 => x"4252414d",
          7887 => x"20202020",
          7888 => x"20202825",
          7889 => x"3038583a",
          7890 => x"25303858",
          7891 => x"292e0a00",
          7892 => x"20202020",
          7893 => x"52414d20",
          7894 => x"20202020",
          7895 => x"20202825",
          7896 => x"3038583a",
          7897 => x"25303858",
          7898 => x"292e0a00",
          7899 => x"20202020",
          7900 => x"53442043",
          7901 => x"41524420",
          7902 => x"20202844",
          7903 => x"65766963",
          7904 => x"6573203d",
          7905 => x"25303264",
          7906 => x"292e0a00",
          7907 => x"20202020",
          7908 => x"54494d45",
          7909 => x"52312020",
          7910 => x"20202854",
          7911 => x"696d6572",
          7912 => x"7320203d",
          7913 => x"25303264",
          7914 => x"292e0a00",
          7915 => x"20202020",
          7916 => x"494e5452",
          7917 => x"20435452",
          7918 => x"4c202843",
          7919 => x"68616e6e",
          7920 => x"656c733d",
          7921 => x"25303264",
          7922 => x"292e0a00",
          7923 => x"20202020",
          7924 => x"57495348",
          7925 => x"424f4e45",
          7926 => x"20425553",
          7927 => x"0a000000",
          7928 => x"20202020",
          7929 => x"57422049",
          7930 => x"32430a00",
          7931 => x"20202020",
          7932 => x"494f4354",
          7933 => x"4c0a0000",
          7934 => x"20202020",
          7935 => x"5053320a",
          7936 => x"00000000",
          7937 => x"20202020",
          7938 => x"5350490a",
          7939 => x"00000000",
          7940 => x"41646472",
          7941 => x"65737365",
          7942 => x"733a0a00",
          7943 => x"20202020",
          7944 => x"43505520",
          7945 => x"52657365",
          7946 => x"74205665",
          7947 => x"63746f72",
          7948 => x"20416464",
          7949 => x"72657373",
          7950 => x"203d2025",
          7951 => x"3038580a",
          7952 => x"00000000",
          7953 => x"20202020",
          7954 => x"43505520",
          7955 => x"4d656d6f",
          7956 => x"72792053",
          7957 => x"74617274",
          7958 => x"20416464",
          7959 => x"72657373",
          7960 => x"203d2025",
          7961 => x"3038580a",
          7962 => x"00000000",
          7963 => x"20202020",
          7964 => x"53746163",
          7965 => x"6b205374",
          7966 => x"61727420",
          7967 => x"41646472",
          7968 => x"65737320",
          7969 => x"20202020",
          7970 => x"203d2025",
          7971 => x"3038580a",
          7972 => x"00000000",
          7973 => x"4d697363",
          7974 => x"3a0a0000",
          7975 => x"20202020",
          7976 => x"5a505520",
          7977 => x"49642020",
          7978 => x"20202020",
          7979 => x"20202020",
          7980 => x"20202020",
          7981 => x"20202020",
          7982 => x"203d2025",
          7983 => x"3034580a",
          7984 => x"00000000",
          7985 => x"20202020",
          7986 => x"53797374",
          7987 => x"656d2043",
          7988 => x"6c6f636b",
          7989 => x"20467265",
          7990 => x"71202020",
          7991 => x"20202020",
          7992 => x"203d2025",
          7993 => x"642e2530",
          7994 => x"34644d48",
          7995 => x"7a0a0000",
          7996 => x"20202020",
          7997 => x"53445241",
          7998 => x"4d20436c",
          7999 => x"6f636b20",
          8000 => x"46726571",
          8001 => x"20202020",
          8002 => x"20202020",
          8003 => x"203d2025",
          8004 => x"642e2530",
          8005 => x"34644d48",
          8006 => x"7a0a0000",
          8007 => x"20202020",
          8008 => x"57697368",
          8009 => x"626f6e65",
          8010 => x"20534452",
          8011 => x"414d2043",
          8012 => x"6c6f636b",
          8013 => x"20467265",
          8014 => x"713d2025",
          8015 => x"642e2530",
          8016 => x"34644d48",
          8017 => x"7a0a0000",
          8018 => x"536d616c",
          8019 => x"6c000000",
          8020 => x"4d656469",
          8021 => x"756d0000",
          8022 => x"466c6578",
          8023 => x"00000000",
          8024 => x"45564f00",
          8025 => x"45564f6d",
          8026 => x"696e0000",
          8027 => x"556e6b6e",
          8028 => x"6f776e00",
          8029 => x"00007ed0",
          8030 => x"01000000",
          8031 => x"00000002",
          8032 => x"00007ecc",
          8033 => x"01000000",
          8034 => x"00000003",
          8035 => x"00007ec8",
          8036 => x"01000000",
          8037 => x"00000004",
          8038 => x"00007ec4",
          8039 => x"01000000",
          8040 => x"00000005",
          8041 => x"00007ec0",
          8042 => x"01000000",
          8043 => x"00000006",
          8044 => x"00007ebc",
          8045 => x"01000000",
          8046 => x"00000007",
          8047 => x"00007eb8",
          8048 => x"01000000",
          8049 => x"00000001",
          8050 => x"00007eb4",
          8051 => x"01000000",
          8052 => x"00000008",
          8053 => x"00007eb0",
          8054 => x"01000000",
          8055 => x"0000000b",
          8056 => x"00007eac",
          8057 => x"01000000",
          8058 => x"00000009",
          8059 => x"00007ea8",
          8060 => x"01000000",
          8061 => x"0000000a",
          8062 => x"00007ea4",
          8063 => x"04000000",
          8064 => x"0000000d",
          8065 => x"00007ea0",
          8066 => x"04000000",
          8067 => x"0000000c",
          8068 => x"00007e9c",
          8069 => x"04000000",
          8070 => x"0000000e",
          8071 => x"00007e98",
          8072 => x"03000000",
          8073 => x"0000000f",
          8074 => x"00007e94",
          8075 => x"04000000",
          8076 => x"0000000f",
          8077 => x"00007e90",
          8078 => x"04000000",
          8079 => x"00000010",
          8080 => x"00007e8c",
          8081 => x"04000000",
          8082 => x"00000011",
          8083 => x"00007e88",
          8084 => x"03000000",
          8085 => x"00000012",
          8086 => x"00007e84",
          8087 => x"03000000",
          8088 => x"00000013",
          8089 => x"00007e80",
          8090 => x"03000000",
          8091 => x"00000014",
          8092 => x"00007e7c",
          8093 => x"03000000",
          8094 => x"00000015",
          8095 => x"1b5b4400",
          8096 => x"1b5b4300",
          8097 => x"1b5b4200",
          8098 => x"1b5b4100",
          8099 => x"1b5b367e",
          8100 => x"1b5b357e",
          8101 => x"1b5b347e",
          8102 => x"1b304600",
          8103 => x"1b5b337e",
          8104 => x"1b5b327e",
          8105 => x"1b5b317e",
          8106 => x"10000000",
          8107 => x"0e000000",
          8108 => x"0d000000",
          8109 => x"0b000000",
          8110 => x"08000000",
          8111 => x"06000000",
          8112 => x"05000000",
          8113 => x"04000000",
          8114 => x"03000000",
          8115 => x"02000000",
          8116 => x"01000000",
          8117 => x"68697374",
          8118 => x"6f727900",
          8119 => x"68697374",
          8120 => x"00000000",
          8121 => x"21000000",
          8122 => x"25303464",
          8123 => x"20202573",
          8124 => x"0a000000",
          8125 => x"4661696c",
          8126 => x"65642074",
          8127 => x"6f207265",
          8128 => x"73657420",
          8129 => x"74686520",
          8130 => x"68697374",
          8131 => x"6f727920",
          8132 => x"66696c65",
          8133 => x"20746f20",
          8134 => x"454f462e",
          8135 => x"0a000000",
          8136 => x"43616e6e",
          8137 => x"6f74206f",
          8138 => x"70656e2f",
          8139 => x"63726561",
          8140 => x"74652068",
          8141 => x"6973746f",
          8142 => x"72792066",
          8143 => x"696c652c",
          8144 => x"20646973",
          8145 => x"61626c69",
          8146 => x"6e672e0a",
          8147 => x"00000000",
          8148 => x"53440000",
          8149 => x"222a2b2c",
          8150 => x"3a3b3c3d",
          8151 => x"3e3f5b5d",
          8152 => x"7c7f0000",
          8153 => x"46415400",
          8154 => x"46415433",
          8155 => x"32000000",
          8156 => x"ebfe904d",
          8157 => x"53444f53",
          8158 => x"352e3000",
          8159 => x"4e4f204e",
          8160 => x"414d4520",
          8161 => x"20202046",
          8162 => x"41543332",
          8163 => x"20202000",
          8164 => x"4e4f204e",
          8165 => x"414d4520",
          8166 => x"20202046",
          8167 => x"41542020",
          8168 => x"20202000",
          8169 => x"00007f50",
          8170 => x"00000000",
          8171 => x"00000000",
          8172 => x"00000000",
          8173 => x"809a4541",
          8174 => x"8e418f80",
          8175 => x"45454549",
          8176 => x"49498e8f",
          8177 => x"9092924f",
          8178 => x"994f5555",
          8179 => x"59999a9b",
          8180 => x"9c9d9e9f",
          8181 => x"41494f55",
          8182 => x"a5a5a6a7",
          8183 => x"a8a9aaab",
          8184 => x"acadaeaf",
          8185 => x"b0b1b2b3",
          8186 => x"b4b5b6b7",
          8187 => x"b8b9babb",
          8188 => x"bcbdbebf",
          8189 => x"c0c1c2c3",
          8190 => x"c4c5c6c7",
          8191 => x"c8c9cacb",
          8192 => x"cccdcecf",
          8193 => x"d0d1d2d3",
          8194 => x"d4d5d6d7",
          8195 => x"d8d9dadb",
          8196 => x"dcdddedf",
          8197 => x"e0e1e2e3",
          8198 => x"e4e5e6e7",
          8199 => x"e8e9eaeb",
          8200 => x"ecedeeef",
          8201 => x"f0f1f2f3",
          8202 => x"f4f5f6f7",
          8203 => x"f8f9fafb",
          8204 => x"fcfdfeff",
          8205 => x"2b2e2c3b",
          8206 => x"3d5b5d2f",
          8207 => x"5c222a3a",
          8208 => x"3c3e3f7c",
          8209 => x"7f000000",
          8210 => x"00010004",
          8211 => x"00100040",
          8212 => x"01000200",
          8213 => x"00000000",
          8214 => x"00010002",
          8215 => x"00040008",
          8216 => x"00100020",
          8217 => x"00000000",
          8218 => x"00000000",
          8219 => x"000074c8",
          8220 => x"01020100",
          8221 => x"00000000",
          8222 => x"00000000",
          8223 => x"000074d0",
          8224 => x"01040100",
          8225 => x"00000000",
          8226 => x"00000000",
          8227 => x"000074d8",
          8228 => x"01140300",
          8229 => x"00000000",
          8230 => x"00000000",
          8231 => x"000074e0",
          8232 => x"012b0300",
          8233 => x"00000000",
          8234 => x"00000000",
          8235 => x"000074e8",
          8236 => x"01300300",
          8237 => x"00000000",
          8238 => x"00000000",
          8239 => x"000074f0",
          8240 => x"013c0400",
          8241 => x"00000000",
          8242 => x"00000000",
          8243 => x"000074f8",
          8244 => x"013d0400",
          8245 => x"00000000",
          8246 => x"00000000",
          8247 => x"00007500",
          8248 => x"013f0400",
          8249 => x"00000000",
          8250 => x"00000000",
          8251 => x"00007508",
          8252 => x"01400400",
          8253 => x"00000000",
          8254 => x"00000000",
          8255 => x"00007510",
          8256 => x"01410400",
          8257 => x"00000000",
          8258 => x"00000000",
          8259 => x"00007514",
          8260 => x"01420400",
          8261 => x"00000000",
          8262 => x"00000000",
          8263 => x"00007518",
          8264 => x"01430400",
          8265 => x"00000000",
          8266 => x"00000000",
          8267 => x"0000751c",
          8268 => x"01500500",
          8269 => x"00000000",
          8270 => x"00000000",
          8271 => x"00007520",
          8272 => x"01510500",
          8273 => x"00000000",
          8274 => x"00000000",
          8275 => x"00007524",
          8276 => x"01540500",
          8277 => x"00000000",
          8278 => x"00000000",
          8279 => x"00007528",
          8280 => x"01550500",
          8281 => x"00000000",
          8282 => x"00000000",
          8283 => x"0000752c",
          8284 => x"01790700",
          8285 => x"00000000",
          8286 => x"00000000",
          8287 => x"00007534",
          8288 => x"01780700",
          8289 => x"00000000",
          8290 => x"00000000",
          8291 => x"00007538",
          8292 => x"01820800",
          8293 => x"00000000",
          8294 => x"00000000",
          8295 => x"00007540",
          8296 => x"01830800",
          8297 => x"00000000",
          8298 => x"00000000",
          8299 => x"00007548",
          8300 => x"01850800",
          8301 => x"00000000",
          8302 => x"00000000",
          8303 => x"00007550",
          8304 => x"01870800",
          8305 => x"00000000",
          8306 => x"00000000",
          8307 => x"00007558",
          8308 => x"018c0900",
          8309 => x"00000000",
          8310 => x"00000000",
          8311 => x"00007560",
          8312 => x"018d0900",
          8313 => x"00000000",
          8314 => x"00000000",
          8315 => x"00007568",
          8316 => x"018e0900",
          8317 => x"00000000",
          8318 => x"00000000",
          8319 => x"00007570",
          8320 => x"018f0900",
          8321 => x"00000000",
          8322 => x"00000000",
          8323 => x"00000000",
          8324 => x"00000000",
          8325 => x"00007fff",
          8326 => x"00000000",
          8327 => x"00007fff",
          8328 => x"00010000",
          8329 => x"00007fff",
          8330 => x"00010000",
          8331 => x"00810000",
          8332 => x"01000000",
          8333 => x"017fffff",
          8334 => x"00000000",
          8335 => x"00000000",
          8336 => x"00007800",
          8337 => x"00000000",
          8338 => x"05f5e100",
          8339 => x"05f5e100",
          8340 => x"05f5e100",
          8341 => x"00000000",
          8342 => x"01010101",
          8343 => x"01010101",
          8344 => x"01011001",
          8345 => x"01000000",
          8346 => x"00000000",
          8347 => x"00000000",
          8348 => x"00000000",
          8349 => x"00000000",
          8350 => x"00000000",
          8351 => x"00000000",
          8352 => x"00000000",
          8353 => x"00000000",
          8354 => x"00000000",
          8355 => x"00000000",
          8356 => x"00000000",
          8357 => x"00000000",
          8358 => x"00000000",
          8359 => x"00000000",
          8360 => x"00000000",
          8361 => x"00000000",
          8362 => x"00000000",
          8363 => x"00000000",
          8364 => x"00000000",
          8365 => x"00000000",
          8366 => x"00000000",
          8367 => x"00000000",
          8368 => x"00000000",
          8369 => x"00000000",
          8370 => x"00007ed4",
          8371 => x"01000000",
          8372 => x"00007edc",
          8373 => x"01000000",
          8374 => x"00007ee4",
          8375 => x"02000000",
          8376 => x"00000000",
          8377 => x"00000000",
          8378 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

