-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b83ff",
          2049 => x"f80d0b0b",
          2050 => x"0b939b04",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b92",
          2121 => x"ff040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b92e2",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b81e7",
          2210 => x"fc738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"92e70400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0b99",
          2219 => x"fb2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0b9b",
          2227 => x"e72d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"95040b0b",
          2317 => x"0b8ca504",
          2318 => x"0b0b0b8c",
          2319 => x"b5040b0b",
          2320 => x"0b8cc504",
          2321 => x"0b0b0b8c",
          2322 => x"d5040b0b",
          2323 => x"0b8ce504",
          2324 => x"0b0b0b8c",
          2325 => x"f5040b0b",
          2326 => x"0b8d8504",
          2327 => x"0b0b0b8d",
          2328 => x"95040b0b",
          2329 => x"0b8da504",
          2330 => x"0b0b0b8d",
          2331 => x"b5040b0b",
          2332 => x"0b8dc504",
          2333 => x"0b0b0b8d",
          2334 => x"d5040b0b",
          2335 => x"0b8de504",
          2336 => x"0b0b0b8d",
          2337 => x"f5040b0b",
          2338 => x"0b8e8404",
          2339 => x"0b0b0b8e",
          2340 => x"93040b0b",
          2341 => x"0b8ea204",
          2342 => x"0b0b0b8e",
          2343 => x"b2040b0b",
          2344 => x"0b8ec204",
          2345 => x"0b0b0b8e",
          2346 => x"d2040b0b",
          2347 => x"0b8ee204",
          2348 => x"0b0b0b8e",
          2349 => x"f2040b0b",
          2350 => x"0b8f8204",
          2351 => x"0b0b0b8f",
          2352 => x"92040b0b",
          2353 => x"0b8fa204",
          2354 => x"0b0b0b8f",
          2355 => x"b2040b0b",
          2356 => x"0b8fc204",
          2357 => x"0b0b0b8f",
          2358 => x"d2040b0b",
          2359 => x"0b8fe204",
          2360 => x"0b0b0b8f",
          2361 => x"f2040b0b",
          2362 => x"0b908204",
          2363 => x"0b0b0b90",
          2364 => x"92040b0b",
          2365 => x"0b90a204",
          2366 => x"0b0b0b90",
          2367 => x"b2040b0b",
          2368 => x"0b90c204",
          2369 => x"0b0b0b90",
          2370 => x"d2040b0b",
          2371 => x"0b90e204",
          2372 => x"0b0b0b90",
          2373 => x"f2040b0b",
          2374 => x"0b918204",
          2375 => x"0b0b0b91",
          2376 => x"92040b0b",
          2377 => x"0b91a204",
          2378 => x"0b0b0b91",
          2379 => x"b2040b0b",
          2380 => x"0b91c204",
          2381 => x"0b0b0b91",
          2382 => x"d2040b0b",
          2383 => x"0b91e204",
          2384 => x"0b0b0b91",
          2385 => x"f2040b0b",
          2386 => x"0b928204",
          2387 => x"0b0b0b92",
          2388 => x"91040b0b",
          2389 => x"0b92a004",
          2390 => x"0b0b0b92",
          2391 => x"b004ffff",
          2392 => x"ffffffff",
          2393 => x"ffffffff",
          2394 => x"ffffffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"048285f8",
          2434 => x"0c80c18c",
          2435 => x"2d8285f8",
          2436 => x"0882a090",
          2437 => x"048285f8",
          2438 => x"0c80ce8e",
          2439 => x"2d8285f8",
          2440 => x"0882a090",
          2441 => x"048285f8",
          2442 => x"0c80cecd",
          2443 => x"2d8285f8",
          2444 => x"0882a090",
          2445 => x"048285f8",
          2446 => x"0c80ceeb",
          2447 => x"2d8285f8",
          2448 => x"0882a090",
          2449 => x"048285f8",
          2450 => x"0c80d5b5",
          2451 => x"2d8285f8",
          2452 => x"0882a090",
          2453 => x"048285f8",
          2454 => x"0c80d6b6",
          2455 => x"2d8285f8",
          2456 => x"0882a090",
          2457 => x"048285f8",
          2458 => x"0c80cf8e",
          2459 => x"2d8285f8",
          2460 => x"0882a090",
          2461 => x"048285f8",
          2462 => x"0c80d6d3",
          2463 => x"2d8285f8",
          2464 => x"0882a090",
          2465 => x"048285f8",
          2466 => x"0c80d8cf",
          2467 => x"2d8285f8",
          2468 => x"0882a090",
          2469 => x"048285f8",
          2470 => x"0c80d4db",
          2471 => x"2d8285f8",
          2472 => x"0882a090",
          2473 => x"048285f8",
          2474 => x"0c80cfc0",
          2475 => x"2d8285f8",
          2476 => x"0882a090",
          2477 => x"048285f8",
          2478 => x"0c80d4f1",
          2479 => x"2d8285f8",
          2480 => x"0882a090",
          2481 => x"048285f8",
          2482 => x"0c80d595",
          2483 => x"2d8285f8",
          2484 => x"0882a090",
          2485 => x"048285f8",
          2486 => x"0c80c395",
          2487 => x"2d8285f8",
          2488 => x"0882a090",
          2489 => x"048285f8",
          2490 => x"0c80c3e4",
          2491 => x"2d8285f8",
          2492 => x"0882a090",
          2493 => x"048285f8",
          2494 => x"0cbbc42d",
          2495 => x"8285f808",
          2496 => x"82a09004",
          2497 => x"8285f80c",
          2498 => x"bdbd2d82",
          2499 => x"85f80882",
          2500 => x"a0900482",
          2501 => x"85f80cbe",
          2502 => x"f02d8285",
          2503 => x"f80882a0",
          2504 => x"90048285",
          2505 => x"f80c81aa",
          2506 => x"bc2d8285",
          2507 => x"f80882a0",
          2508 => x"90048285",
          2509 => x"f80c81b7",
          2510 => x"af2d8285",
          2511 => x"f80882a0",
          2512 => x"90048285",
          2513 => x"f80c81af",
          2514 => x"a32d8285",
          2515 => x"f80882a0",
          2516 => x"90048285",
          2517 => x"f80c81b2",
          2518 => x"a02d8285",
          2519 => x"f80882a0",
          2520 => x"90048285",
          2521 => x"f80c81bc",
          2522 => x"bd2d8285",
          2523 => x"f80882a0",
          2524 => x"90048285",
          2525 => x"f80c81c5",
          2526 => x"a82d8285",
          2527 => x"f80882a0",
          2528 => x"90048285",
          2529 => x"f80c81b6",
          2530 => x"912d8285",
          2531 => x"f80882a0",
          2532 => x"90048285",
          2533 => x"f80c81bf",
          2534 => x"de2d8285",
          2535 => x"f80882a0",
          2536 => x"90048285",
          2537 => x"f80c81c0",
          2538 => x"fd2d8285",
          2539 => x"f80882a0",
          2540 => x"90048285",
          2541 => x"f80c81c1",
          2542 => x"9c2d8285",
          2543 => x"f80882a0",
          2544 => x"90048285",
          2545 => x"f80c81c9",
          2546 => x"912d8285",
          2547 => x"f80882a0",
          2548 => x"90048285",
          2549 => x"f80c81c6",
          2550 => x"f52d8285",
          2551 => x"f80882a0",
          2552 => x"90048285",
          2553 => x"f80c81cb",
          2554 => x"e52d8285",
          2555 => x"f80882a0",
          2556 => x"90048285",
          2557 => x"f80c81c2",
          2558 => x"a22d8285",
          2559 => x"f80882a0",
          2560 => x"90048285",
          2561 => x"f80c81ce",
          2562 => x"e52d8285",
          2563 => x"f80882a0",
          2564 => x"90048285",
          2565 => x"f80c81cf",
          2566 => x"e62d8285",
          2567 => x"f80882a0",
          2568 => x"90048285",
          2569 => x"f80c81b8",
          2570 => x"8f2d8285",
          2571 => x"f80882a0",
          2572 => x"90048285",
          2573 => x"f80c81b7",
          2574 => x"e82d8285",
          2575 => x"f80882a0",
          2576 => x"90048285",
          2577 => x"f80c81b9",
          2578 => x"932d8285",
          2579 => x"f80882a0",
          2580 => x"90048285",
          2581 => x"f80c81c2",
          2582 => x"f92d8285",
          2583 => x"f80882a0",
          2584 => x"90048285",
          2585 => x"f80c81d0",
          2586 => x"d72d8285",
          2587 => x"f80882a0",
          2588 => x"90048285",
          2589 => x"f80c81d2",
          2590 => x"e52d8285",
          2591 => x"f80882a0",
          2592 => x"90048285",
          2593 => x"f80c81d6",
          2594 => x"a72d8285",
          2595 => x"f80882a0",
          2596 => x"90048285",
          2597 => x"f80c81a9",
          2598 => x"db2d8285",
          2599 => x"f80882a0",
          2600 => x"90048285",
          2601 => x"f80c81d9",
          2602 => x"952d8285",
          2603 => x"f80882a0",
          2604 => x"90048285",
          2605 => x"f80c81e7",
          2606 => x"d92d8285",
          2607 => x"f80882a0",
          2608 => x"90048285",
          2609 => x"f80c81e5",
          2610 => x"c02d8285",
          2611 => x"f80882a0",
          2612 => x"90048285",
          2613 => x"f80c80fa",
          2614 => x"e82d8285",
          2615 => x"f80882a0",
          2616 => x"90048285",
          2617 => x"f80c80fc",
          2618 => x"d22d8285",
          2619 => x"f80882a0",
          2620 => x"90048285",
          2621 => x"f80c80fe",
          2622 => x"b62d8285",
          2623 => x"f80882a0",
          2624 => x"90048285",
          2625 => x"f80cbbed",
          2626 => x"2d8285f8",
          2627 => x"0882a090",
          2628 => x"048285f8",
          2629 => x"0cbd932d",
          2630 => x"8285f808",
          2631 => x"82a09004",
          2632 => x"8285f80c",
          2633 => x"80c0802d",
          2634 => x"8285f808",
          2635 => x"82a09004",
          2636 => x"8285f80c",
          2637 => x"a1fd2d82",
          2638 => x"85f80882",
          2639 => x"a090043c",
          2640 => x"04000010",
          2641 => x"10101010",
          2642 => x"10101010",
          2643 => x"10101010",
          2644 => x"10101010",
          2645 => x"10101010",
          2646 => x"10101010",
          2647 => x"10101010",
          2648 => x"10105351",
          2649 => x"04000073",
          2650 => x"81ff0673",
          2651 => x"83060981",
          2652 => x"05830510",
          2653 => x"10102b07",
          2654 => x"72fc060c",
          2655 => x"51510472",
          2656 => x"72807281",
          2657 => x"06ff0509",
          2658 => x"72060571",
          2659 => x"1052720a",
          2660 => x"100a5372",
          2661 => x"ed385151",
          2662 => x"53510482",
          2663 => x"85ec7082",
          2664 => x"9da8278e",
          2665 => x"38807170",
          2666 => x"8405530c",
          2667 => x"0b0b0b93",
          2668 => x"9e048c81",
          2669 => x"51ba9d04",
          2670 => x"008285f8",
          2671 => x"08028285",
          2672 => x"f80cfe3d",
          2673 => x"0d8285f8",
          2674 => x"08880508",
          2675 => x"8285f808",
          2676 => x"fc050c82",
          2677 => x"85f808fc",
          2678 => x"05085271",
          2679 => x"338285f8",
          2680 => x"08fc0508",
          2681 => x"81058285",
          2682 => x"f808fc05",
          2683 => x"0c7081ff",
          2684 => x"06515170",
          2685 => x"802e8338",
          2686 => x"da398285",
          2687 => x"f808fc05",
          2688 => x"08ff0582",
          2689 => x"85f808fc",
          2690 => x"050c8285",
          2691 => x"f808fc05",
          2692 => x"088285f8",
          2693 => x"08880508",
          2694 => x"31708285",
          2695 => x"ec0c5184",
          2696 => x"3d0d8285",
          2697 => x"f80c0482",
          2698 => x"85f80802",
          2699 => x"8285f80c",
          2700 => x"fe3d0d82",
          2701 => x"85f80888",
          2702 => x"05088285",
          2703 => x"f808fc05",
          2704 => x"0c8285f8",
          2705 => x"088c0508",
          2706 => x"52713382",
          2707 => x"85f8088c",
          2708 => x"05088105",
          2709 => x"8285f808",
          2710 => x"8c050c82",
          2711 => x"85f808fc",
          2712 => x"05085351",
          2713 => x"70723482",
          2714 => x"85f808fc",
          2715 => x"05088105",
          2716 => x"8285f808",
          2717 => x"fc050c70",
          2718 => x"81ff0651",
          2719 => x"70802e84",
          2720 => x"38ffbe39",
          2721 => x"8285f808",
          2722 => x"88050870",
          2723 => x"8285ec0c",
          2724 => x"51843d0d",
          2725 => x"8285f80c",
          2726 => x"048285f8",
          2727 => x"08028285",
          2728 => x"f80cfd3d",
          2729 => x"0d8285f8",
          2730 => x"08880508",
          2731 => x"8285f808",
          2732 => x"fc050c82",
          2733 => x"85f8088c",
          2734 => x"05088285",
          2735 => x"f808f805",
          2736 => x"0c8285f8",
          2737 => x"08900508",
          2738 => x"802e80e5",
          2739 => x"388285f8",
          2740 => x"08900508",
          2741 => x"81058285",
          2742 => x"f8089005",
          2743 => x"0c8285f8",
          2744 => x"08900508",
          2745 => x"ff058285",
          2746 => x"f8089005",
          2747 => x"0c8285f8",
          2748 => x"08900508",
          2749 => x"802eba38",
          2750 => x"8285f808",
          2751 => x"f8050851",
          2752 => x"70338285",
          2753 => x"f808f805",
          2754 => x"08810582",
          2755 => x"85f808f8",
          2756 => x"050c8285",
          2757 => x"f808fc05",
          2758 => x"08525271",
          2759 => x"71348285",
          2760 => x"f808fc05",
          2761 => x"08810582",
          2762 => x"85f808fc",
          2763 => x"050cffad",
          2764 => x"398285f8",
          2765 => x"08880508",
          2766 => x"708285ec",
          2767 => x"0c51853d",
          2768 => x"0d8285f8",
          2769 => x"0c048285",
          2770 => x"f8080282",
          2771 => x"85f80cfd",
          2772 => x"3d0d8285",
          2773 => x"f8089005",
          2774 => x"08802e81",
          2775 => x"f4388285",
          2776 => x"f8088c05",
          2777 => x"08527133",
          2778 => x"8285f808",
          2779 => x"8c050881",
          2780 => x"058285f8",
          2781 => x"088c050c",
          2782 => x"8285f808",
          2783 => x"88050870",
          2784 => x"337281ff",
          2785 => x"06535454",
          2786 => x"5171712e",
          2787 => x"843880ce",
          2788 => x"398285f8",
          2789 => x"08880508",
          2790 => x"52713382",
          2791 => x"85f80888",
          2792 => x"05088105",
          2793 => x"8285f808",
          2794 => x"88050c70",
          2795 => x"81ff0651",
          2796 => x"51708d38",
          2797 => x"800b8285",
          2798 => x"f808fc05",
          2799 => x"0c819b39",
          2800 => x"8285f808",
          2801 => x"900508ff",
          2802 => x"058285f8",
          2803 => x"0890050c",
          2804 => x"8285f808",
          2805 => x"90050880",
          2806 => x"2e8438ff",
          2807 => x"81398285",
          2808 => x"f8089005",
          2809 => x"08802e80",
          2810 => x"e8388285",
          2811 => x"f8088805",
          2812 => x"08703352",
          2813 => x"53708d38",
          2814 => x"ff0b8285",
          2815 => x"f808fc05",
          2816 => x"0c80d739",
          2817 => x"8285f808",
          2818 => x"8c0508ff",
          2819 => x"058285f8",
          2820 => x"088c050c",
          2821 => x"8285f808",
          2822 => x"8c050870",
          2823 => x"33525270",
          2824 => x"8c38810b",
          2825 => x"8285f808",
          2826 => x"fc050cae",
          2827 => x"398285f8",
          2828 => x"08880508",
          2829 => x"70338285",
          2830 => x"f8088c05",
          2831 => x"08703372",
          2832 => x"71317082",
          2833 => x"85f808fc",
          2834 => x"050c5355",
          2835 => x"5252538a",
          2836 => x"39800b82",
          2837 => x"85f808fc",
          2838 => x"050c8285",
          2839 => x"f808fc05",
          2840 => x"088285ec",
          2841 => x"0c853d0d",
          2842 => x"8285f80c",
          2843 => x"048285f8",
          2844 => x"08028285",
          2845 => x"f80cfe3d",
          2846 => x"0d8285f8",
          2847 => x"08880508",
          2848 => x"8285f808",
          2849 => x"fc050c82",
          2850 => x"85f80890",
          2851 => x"0508802e",
          2852 => x"80d43882",
          2853 => x"85f80890",
          2854 => x"05088105",
          2855 => x"8285f808",
          2856 => x"90050c82",
          2857 => x"85f80890",
          2858 => x"0508ff05",
          2859 => x"8285f808",
          2860 => x"90050c82",
          2861 => x"85f80890",
          2862 => x"0508802e",
          2863 => x"a9388285",
          2864 => x"f8088c05",
          2865 => x"08517082",
          2866 => x"85f808fc",
          2867 => x"05085252",
          2868 => x"71713482",
          2869 => x"85f808fc",
          2870 => x"05088105",
          2871 => x"8285f808",
          2872 => x"fc050cff",
          2873 => x"be398285",
          2874 => x"f8088805",
          2875 => x"08708285",
          2876 => x"ec0c5184",
          2877 => x"3d0d8285",
          2878 => x"f80c0482",
          2879 => x"85f80802",
          2880 => x"8285f80c",
          2881 => x"f93d0d80",
          2882 => x"0b8285f8",
          2883 => x"08fc050c",
          2884 => x"8285f808",
          2885 => x"88050880",
          2886 => x"25b93882",
          2887 => x"85f80888",
          2888 => x"05083082",
          2889 => x"85f80888",
          2890 => x"050c800b",
          2891 => x"8285f808",
          2892 => x"f4050c82",
          2893 => x"85f808fc",
          2894 => x"05088a38",
          2895 => x"810b8285",
          2896 => x"f808f405",
          2897 => x"0c8285f8",
          2898 => x"08f40508",
          2899 => x"8285f808",
          2900 => x"fc050c82",
          2901 => x"85f8088c",
          2902 => x"05088025",
          2903 => x"b9388285",
          2904 => x"f8088c05",
          2905 => x"08308285",
          2906 => x"f8088c05",
          2907 => x"0c800b82",
          2908 => x"85f808f0",
          2909 => x"050c8285",
          2910 => x"f808fc05",
          2911 => x"088a3881",
          2912 => x"0b8285f8",
          2913 => x"08f0050c",
          2914 => x"8285f808",
          2915 => x"f0050882",
          2916 => x"85f808fc",
          2917 => x"050c8053",
          2918 => x"8285f808",
          2919 => x"8c050852",
          2920 => x"8285f808",
          2921 => x"88050851",
          2922 => x"83c53f82",
          2923 => x"85ec0870",
          2924 => x"8285f808",
          2925 => x"f8050c54",
          2926 => x"8285f808",
          2927 => x"fc050880",
          2928 => x"2e903882",
          2929 => x"85f808f8",
          2930 => x"05083082",
          2931 => x"85f808f8",
          2932 => x"050c8285",
          2933 => x"f808f805",
          2934 => x"08708285",
          2935 => x"ec0c5489",
          2936 => x"3d0d8285",
          2937 => x"f80c0482",
          2938 => x"85f80802",
          2939 => x"8285f80c",
          2940 => x"fb3d0d80",
          2941 => x"0b8285f8",
          2942 => x"08fc050c",
          2943 => x"8285f808",
          2944 => x"88050880",
          2945 => x"25993882",
          2946 => x"85f80888",
          2947 => x"05083082",
          2948 => x"85f80888",
          2949 => x"050c810b",
          2950 => x"8285f808",
          2951 => x"fc050c82",
          2952 => x"85f8088c",
          2953 => x"05088025",
          2954 => x"90388285",
          2955 => x"f8088c05",
          2956 => x"08308285",
          2957 => x"f8088c05",
          2958 => x"0c815382",
          2959 => x"85f8088c",
          2960 => x"05085282",
          2961 => x"85f80888",
          2962 => x"05085182",
          2963 => x"a23f8285",
          2964 => x"ec087082",
          2965 => x"85f808f8",
          2966 => x"050c5482",
          2967 => x"85f808fc",
          2968 => x"0508802e",
          2969 => x"90388285",
          2970 => x"f808f805",
          2971 => x"08308285",
          2972 => x"f808f805",
          2973 => x"0c8285f8",
          2974 => x"08f80508",
          2975 => x"708285ec",
          2976 => x"0c54873d",
          2977 => x"0d8285f8",
          2978 => x"0c048285",
          2979 => x"f8080282",
          2980 => x"85f80cff",
          2981 => x"3d0d800b",
          2982 => x"8285f808",
          2983 => x"fc050c82",
          2984 => x"85f80888",
          2985 => x"05088106",
          2986 => x"ff117009",
          2987 => x"708285f8",
          2988 => x"088c0508",
          2989 => x"068285f8",
          2990 => x"08fc0508",
          2991 => x"118285f8",
          2992 => x"08fc050c",
          2993 => x"8285f808",
          2994 => x"88050881",
          2995 => x"2a8285f8",
          2996 => x"0888050c",
          2997 => x"8285f808",
          2998 => x"8c050810",
          2999 => x"8285f808",
          3000 => x"8c050c51",
          3001 => x"51515182",
          3002 => x"85f80888",
          3003 => x"0508802e",
          3004 => x"8438ffab",
          3005 => x"398285f8",
          3006 => x"08fc0508",
          3007 => x"708285ec",
          3008 => x"0c51833d",
          3009 => x"0d8285f8",
          3010 => x"0c048285",
          3011 => x"f8080282",
          3012 => x"85f80cfd",
          3013 => x"3d0d8053",
          3014 => x"8285f808",
          3015 => x"8c050852",
          3016 => x"8285f808",
          3017 => x"88050851",
          3018 => x"80c53f82",
          3019 => x"85ec0870",
          3020 => x"8285ec0c",
          3021 => x"54853d0d",
          3022 => x"8285f80c",
          3023 => x"048285f8",
          3024 => x"08028285",
          3025 => x"f80cfd3d",
          3026 => x"0d815382",
          3027 => x"85f8088c",
          3028 => x"05085282",
          3029 => x"85f80888",
          3030 => x"05085193",
          3031 => x"3f8285ec",
          3032 => x"08708285",
          3033 => x"ec0c5485",
          3034 => x"3d0d8285",
          3035 => x"f80c0482",
          3036 => x"85f80802",
          3037 => x"8285f80c",
          3038 => x"fd3d0d81",
          3039 => x"0b8285f8",
          3040 => x"08fc050c",
          3041 => x"800b8285",
          3042 => x"f808f805",
          3043 => x"0c8285f8",
          3044 => x"088c0508",
          3045 => x"8285f808",
          3046 => x"88050827",
          3047 => x"b9388285",
          3048 => x"f808fc05",
          3049 => x"08802eae",
          3050 => x"38800b82",
          3051 => x"85f8088c",
          3052 => x"050824a2",
          3053 => x"388285f8",
          3054 => x"088c0508",
          3055 => x"108285f8",
          3056 => x"088c050c",
          3057 => x"8285f808",
          3058 => x"fc050810",
          3059 => x"8285f808",
          3060 => x"fc050cff",
          3061 => x"b8398285",
          3062 => x"f808fc05",
          3063 => x"08802e80",
          3064 => x"e1388285",
          3065 => x"f8088c05",
          3066 => x"088285f8",
          3067 => x"08880508",
          3068 => x"26ad3882",
          3069 => x"85f80888",
          3070 => x"05088285",
          3071 => x"f8088c05",
          3072 => x"08318285",
          3073 => x"f8088805",
          3074 => x"0c8285f8",
          3075 => x"08f80508",
          3076 => x"8285f808",
          3077 => x"fc050807",
          3078 => x"8285f808",
          3079 => x"f8050c82",
          3080 => x"85f808fc",
          3081 => x"0508812a",
          3082 => x"8285f808",
          3083 => x"fc050c82",
          3084 => x"85f8088c",
          3085 => x"0508812a",
          3086 => x"8285f808",
          3087 => x"8c050cff",
          3088 => x"95398285",
          3089 => x"f8089005",
          3090 => x"08802e93",
          3091 => x"388285f8",
          3092 => x"08880508",
          3093 => x"708285f8",
          3094 => x"08f4050c",
          3095 => x"51913982",
          3096 => x"85f808f8",
          3097 => x"05087082",
          3098 => x"85f808f4",
          3099 => x"050c5182",
          3100 => x"85f808f4",
          3101 => x"05088285",
          3102 => x"ec0c853d",
          3103 => x"0d8285f8",
          3104 => x"0c04f93d",
          3105 => x"0d797008",
          3106 => x"70565658",
          3107 => x"74802e80",
          3108 => x"e3389539",
          3109 => x"750851f2",
          3110 => x"a03f8285",
          3111 => x"ec081578",
          3112 => x"0c851633",
          3113 => x"5480cd39",
          3114 => x"74335473",
          3115 => x"a02e0981",
          3116 => x"06863881",
          3117 => x"1555f139",
          3118 => x"80577684",
          3119 => x"2b8280ec",
          3120 => x"05700852",
          3121 => x"56f1f23f",
          3122 => x"8285ec08",
          3123 => x"53745275",
          3124 => x"0851f4f2",
          3125 => x"3f8285ec",
          3126 => x"088b3884",
          3127 => x"16335473",
          3128 => x"812effb0",
          3129 => x"38811770",
          3130 => x"81ff0658",
          3131 => x"54997727",
          3132 => x"c938ff54",
          3133 => x"738285ec",
          3134 => x"0c893d0d",
          3135 => x"04ff3d0d",
          3136 => x"73527193",
          3137 => x"26818d38",
          3138 => x"71822b52",
          3139 => x"81e88c12",
          3140 => x"080481ea",
          3141 => x"f4518180",
          3142 => x"3981eb80",
          3143 => x"5180f939",
          3144 => x"81eb9451",
          3145 => x"80f23981",
          3146 => x"eba85180",
          3147 => x"eb3981eb",
          3148 => x"b85180e4",
          3149 => x"3981ebc8",
          3150 => x"5180dd39",
          3151 => x"81ebdc51",
          3152 => x"80d63981",
          3153 => x"ebec5180",
          3154 => x"cf3981ec",
          3155 => x"845180c8",
          3156 => x"3981ec9c",
          3157 => x"5180c139",
          3158 => x"81ecb451",
          3159 => x"bb3981ec",
          3160 => x"d051b539",
          3161 => x"81ece451",
          3162 => x"af3981ed",
          3163 => x"9051a939",
          3164 => x"81eda451",
          3165 => x"a33981ed",
          3166 => x"c4519d39",
          3167 => x"81edd851",
          3168 => x"973981ed",
          3169 => x"f0519139",
          3170 => x"81ee8851",
          3171 => x"8b3981ee",
          3172 => x"a0518539",
          3173 => x"81eeac51",
          3174 => x"abd13f83",
          3175 => x"3d0d04fb",
          3176 => x"3d0d7779",
          3177 => x"56567487",
          3178 => x"e7269238",
          3179 => x"87e85275",
          3180 => x"51f9d73f",
          3181 => x"74528285",
          3182 => x"ec085190",
          3183 => x"3987e852",
          3184 => x"7451fac6",
          3185 => x"3f8285ec",
          3186 => x"08527551",
          3187 => x"fabc3f82",
          3188 => x"85ec0854",
          3189 => x"79537552",
          3190 => x"81eebc51",
          3191 => x"b0fd3f87",
          3192 => x"3d0d04ec",
          3193 => x"3d0d6602",
          3194 => x"840580e3",
          3195 => x"05335b57",
          3196 => x"80687809",
          3197 => x"8105707a",
          3198 => x"07732551",
          3199 => x"57595978",
          3200 => x"567787ff",
          3201 => x"26833881",
          3202 => x"56747607",
          3203 => x"7081ff06",
          3204 => x"51559356",
          3205 => x"74818638",
          3206 => x"81537652",
          3207 => x"8c3d7052",
          3208 => x"56818698",
          3209 => x"3f8285ec",
          3210 => x"08578285",
          3211 => x"ec08b938",
          3212 => x"8285ec08",
          3213 => x"87c09888",
          3214 => x"0c8285ec",
          3215 => x"0859963d",
          3216 => x"d4055484",
          3217 => x"80537752",
          3218 => x"7551818a",
          3219 => x"d63f8285",
          3220 => x"ec085782",
          3221 => x"85ec0890",
          3222 => x"387a5574",
          3223 => x"802e8938",
          3224 => x"74197519",
          3225 => x"5959d739",
          3226 => x"963dd805",
          3227 => x"518192bf",
          3228 => x"3f760981",
          3229 => x"05707807",
          3230 => x"80257b09",
          3231 => x"8105709f",
          3232 => x"2a720651",
          3233 => x"57515674",
          3234 => x"802e9038",
          3235 => x"81eee053",
          3236 => x"87c09888",
          3237 => x"08527851",
          3238 => x"fe853f76",
          3239 => x"56758285",
          3240 => x"ec0c963d",
          3241 => x"0d04f93d",
          3242 => x"0d7b0284",
          3243 => x"05b30533",
          3244 => x"5758ff57",
          3245 => x"80537a52",
          3246 => x"7951fea7",
          3247 => x"3f8285ec",
          3248 => x"08a43875",
          3249 => x"802e8838",
          3250 => x"75812e98",
          3251 => x"38983960",
          3252 => x"557f5482",
          3253 => x"85ec537e",
          3254 => x"527d5177",
          3255 => x"2d8285ec",
          3256 => x"08578339",
          3257 => x"77047682",
          3258 => x"85ec0c89",
          3259 => x"3d0d04f3",
          3260 => x"3d0d7f61",
          3261 => x"63028c05",
          3262 => x"80cf0533",
          3263 => x"73731568",
          3264 => x"415f5c5c",
          3265 => x"5e5e5e7a",
          3266 => x"5281eee8",
          3267 => x"51aecc3f",
          3268 => x"81eef051",
          3269 => x"a8d53f80",
          3270 => x"55747927",
          3271 => x"80f4387b",
          3272 => x"902e8938",
          3273 => x"7ba02ea4",
          3274 => x"3880c139",
          3275 => x"74185372",
          3276 => x"7a278d38",
          3277 => x"72225281",
          3278 => x"eef451ae",
          3279 => x"9e3f8839",
          3280 => x"81ef8051",
          3281 => x"a8a53f82",
          3282 => x"1555bf39",
          3283 => x"74185372",
          3284 => x"7a278d38",
          3285 => x"72085281",
          3286 => x"eee851ad",
          3287 => x"fe3f8839",
          3288 => x"81eefc51",
          3289 => x"a8853f84",
          3290 => x"15559f39",
          3291 => x"74185372",
          3292 => x"7a278d38",
          3293 => x"72335281",
          3294 => x"ef8851ad",
          3295 => x"de3f8839",
          3296 => x"81ef9051",
          3297 => x"a7e53f81",
          3298 => x"1555a051",
          3299 => x"a7803fff",
          3300 => x"883981ef",
          3301 => x"9451a7d3",
          3302 => x"3f805574",
          3303 => x"7927bb38",
          3304 => x"74187033",
          3305 => x"55538056",
          3306 => x"727a2783",
          3307 => x"38815680",
          3308 => x"539f7427",
          3309 => x"83388153",
          3310 => x"75730670",
          3311 => x"81ff0651",
          3312 => x"5372802e",
          3313 => x"8b387380",
          3314 => x"fe268538",
          3315 => x"73518339",
          3316 => x"a051a6ba",
          3317 => x"3f811555",
          3318 => x"c23981ef",
          3319 => x"9851a78b",
          3320 => x"3f781879",
          3321 => x"1c5c589b",
          3322 => x"fb3f8285",
          3323 => x"ec08982b",
          3324 => x"70982c51",
          3325 => x"5776a02e",
          3326 => x"098106ae",
          3327 => x"389be53f",
          3328 => x"8285ec08",
          3329 => x"982b7098",
          3330 => x"2c70a032",
          3331 => x"70098105",
          3332 => x"729b3270",
          3333 => x"09810570",
          3334 => x"72077375",
          3335 => x"07065158",
          3336 => x"58595751",
          3337 => x"57807324",
          3338 => x"d438769b",
          3339 => x"2e098106",
          3340 => x"85388053",
          3341 => x"8c397c1e",
          3342 => x"53727826",
          3343 => x"fdc938ff",
          3344 => x"53728285",
          3345 => x"ec0c8f3d",
          3346 => x"0d04fc3d",
          3347 => x"0d029b05",
          3348 => x"3381ef9c",
          3349 => x"5381efa0",
          3350 => x"5255abff",
          3351 => x"3f8284c4",
          3352 => x"2251a4d1",
          3353 => x"3f81efac",
          3354 => x"5481efb8",
          3355 => x"538284c5",
          3356 => x"335281ef",
          3357 => x"c051abe3",
          3358 => x"3f74802e",
          3359 => x"8438a086",
          3360 => x"3f863d0d",
          3361 => x"04fe3d0d",
          3362 => x"87c09680",
          3363 => x"0853a4ec",
          3364 => x"3f815196",
          3365 => x"eb3f81ef",
          3366 => x"dc5198e0",
          3367 => x"3f805196",
          3368 => x"df3f7281",
          3369 => x"2a708106",
          3370 => x"51527180",
          3371 => x"2e923881",
          3372 => x"5196cd3f",
          3373 => x"81eff451",
          3374 => x"98c23f80",
          3375 => x"5196c13f",
          3376 => x"72822a70",
          3377 => x"81065152",
          3378 => x"71802e92",
          3379 => x"38815196",
          3380 => x"af3f81f0",
          3381 => x"885198a4",
          3382 => x"3f805196",
          3383 => x"a33f7283",
          3384 => x"2a708106",
          3385 => x"51527180",
          3386 => x"2e923881",
          3387 => x"5196913f",
          3388 => x"81f09851",
          3389 => x"98863f80",
          3390 => x"5196853f",
          3391 => x"72842a70",
          3392 => x"81065152",
          3393 => x"71802e92",
          3394 => x"38815195",
          3395 => x"f33f81f0",
          3396 => x"ac5197e8",
          3397 => x"3f805195",
          3398 => x"e73f7285",
          3399 => x"2a708106",
          3400 => x"51527180",
          3401 => x"2e923881",
          3402 => x"5195d53f",
          3403 => x"81f0c051",
          3404 => x"97ca3f80",
          3405 => x"5195c93f",
          3406 => x"72862a70",
          3407 => x"81065152",
          3408 => x"71802e92",
          3409 => x"38815195",
          3410 => x"b73f81f0",
          3411 => x"d45197ac",
          3412 => x"3f805195",
          3413 => x"ab3f7287",
          3414 => x"2a708106",
          3415 => x"51527180",
          3416 => x"2e923881",
          3417 => x"5195993f",
          3418 => x"81f0e851",
          3419 => x"978e3f80",
          3420 => x"51958d3f",
          3421 => x"72882a70",
          3422 => x"81065152",
          3423 => x"71802e92",
          3424 => x"38815194",
          3425 => x"fb3f81f0",
          3426 => x"fc5196f0",
          3427 => x"3f805194",
          3428 => x"ef3fa2f0",
          3429 => x"3f843d0d",
          3430 => x"04fb3d0d",
          3431 => x"77028405",
          3432 => x"a3053370",
          3433 => x"55565680",
          3434 => x"527551ed",
          3435 => x"c03f0b0b",
          3436 => x"8280e833",
          3437 => x"5473ab38",
          3438 => x"815381f1",
          3439 => x"bc52829c",
          3440 => x"cc5180fe",
          3441 => x"f73f8285",
          3442 => x"ec080981",
          3443 => x"05708285",
          3444 => x"ec080780",
          3445 => x"25827131",
          3446 => x"51515473",
          3447 => x"0b0b8280",
          3448 => x"e8340b0b",
          3449 => x"8280e833",
          3450 => x"5473812e",
          3451 => x"098106af",
          3452 => x"38829ccc",
          3453 => x"53745275",
          3454 => x"5181b9c4",
          3455 => x"3f8285ec",
          3456 => x"08802e8b",
          3457 => x"388285ec",
          3458 => x"0851a2df",
          3459 => x"3f913982",
          3460 => x"9ccc5181",
          3461 => x"8b993f82",
          3462 => x"0b0b0b82",
          3463 => x"80e8340b",
          3464 => x"0b8280e8",
          3465 => x"33547382",
          3466 => x"2e098106",
          3467 => x"8c3881f1",
          3468 => x"cc537452",
          3469 => x"7551b592",
          3470 => x"3f800b82",
          3471 => x"85ec0c87",
          3472 => x"3d0d04ce",
          3473 => x"3d0d8070",
          3474 => x"71829cc8",
          3475 => x"0c5f5d81",
          3476 => x"527c5180",
          3477 => x"cd933f82",
          3478 => x"85ec0881",
          3479 => x"ff065978",
          3480 => x"7d2e0981",
          3481 => x"06a13881",
          3482 => x"f1d45296",
          3483 => x"3d705259",
          3484 => x"a7ff3f7c",
          3485 => x"53785282",
          3486 => x"86f85180",
          3487 => x"fcdd3f82",
          3488 => x"85ec087d",
          3489 => x"2e883881",
          3490 => x"f1d8518d",
          3491 => x"8a398170",
          3492 => x"5f5d81f2",
          3493 => x"9051a1d3",
          3494 => x"3f963d70",
          3495 => x"465a80f8",
          3496 => x"527951fd",
          3497 => x"f43fb43d",
          3498 => x"ff840551",
          3499 => x"f3d43f82",
          3500 => x"85ec0890",
          3501 => x"2b70902c",
          3502 => x"51597880",
          3503 => x"c22e879c",
          3504 => x"387880c2",
          3505 => x"24b23878",
          3506 => x"bd2e81d1",
          3507 => x"3878bd24",
          3508 => x"90387880",
          3509 => x"2effbb38",
          3510 => x"78bc2e80",
          3511 => x"da388abb",
          3512 => x"397880c0",
          3513 => x"2e839438",
          3514 => x"7880c024",
          3515 => x"85cd3878",
          3516 => x"bf2e828a",
          3517 => x"388aa439",
          3518 => x"7880f92e",
          3519 => x"89c33878",
          3520 => x"80f92492",
          3521 => x"387880c3",
          3522 => x"2e87fa38",
          3523 => x"7880f82e",
          3524 => x"898c388a",
          3525 => x"86397881",
          3526 => x"832e89ed",
          3527 => x"38788183",
          3528 => x"248b3878",
          3529 => x"81822e89",
          3530 => x"d33889ef",
          3531 => x"39788185",
          3532 => x"2e89e238",
          3533 => x"89e539b4",
          3534 => x"3dff8011",
          3535 => x"53ff8405",
          3536 => x"51a8903f",
          3537 => x"8285ec08",
          3538 => x"802efec6",
          3539 => x"38b43dfe",
          3540 => x"fc1153ff",
          3541 => x"840551a7",
          3542 => x"fa3f8285",
          3543 => x"ec08802e",
          3544 => x"feb038b4",
          3545 => x"3dfef811",
          3546 => x"53ff8405",
          3547 => x"51a7e43f",
          3548 => x"8285ec08",
          3549 => x"86388285",
          3550 => x"ec084281",
          3551 => x"f294519f",
          3552 => x"ea3f6363",
          3553 => x"5c5a797b",
          3554 => x"2781e938",
          3555 => x"6159787a",
          3556 => x"7084055c",
          3557 => x"0c7a7a26",
          3558 => x"f53881d8",
          3559 => x"39b43dff",
          3560 => x"801153ff",
          3561 => x"840551a7",
          3562 => x"aa3f8285",
          3563 => x"ec08802e",
          3564 => x"fde038b4",
          3565 => x"3dfefc11",
          3566 => x"53ff8405",
          3567 => x"51a7943f",
          3568 => x"8285ec08",
          3569 => x"802efdca",
          3570 => x"38b43dfe",
          3571 => x"f81153ff",
          3572 => x"840551a6",
          3573 => x"fe3f8285",
          3574 => x"ec08802e",
          3575 => x"fdb43881",
          3576 => x"f2a4519f",
          3577 => x"863f635a",
          3578 => x"79632781",
          3579 => x"87386159",
          3580 => x"79708105",
          3581 => x"5b337934",
          3582 => x"61810542",
          3583 => x"eb39b43d",
          3584 => x"ff801153",
          3585 => x"ff840551",
          3586 => x"a6c93f82",
          3587 => x"85ec0880",
          3588 => x"2efcff38",
          3589 => x"b43dfefc",
          3590 => x"1153ff84",
          3591 => x"0551a6b3",
          3592 => x"3f8285ec",
          3593 => x"08802efc",
          3594 => x"e938b43d",
          3595 => x"fef81153",
          3596 => x"ff840551",
          3597 => x"a69d3f82",
          3598 => x"85ec0880",
          3599 => x"2efcd338",
          3600 => x"81f2b051",
          3601 => x"9ea53f63",
          3602 => x"5a796327",
          3603 => x"a7386170",
          3604 => x"337b335e",
          3605 => x"5a5b787c",
          3606 => x"2e913878",
          3607 => x"557a5479",
          3608 => x"33537952",
          3609 => x"81f2c051",
          3610 => x"a3f13f81",
          3611 => x"1a628105",
          3612 => x"435ad639",
          3613 => x"81f2d851",
          3614 => x"82bb39b4",
          3615 => x"3dff8011",
          3616 => x"53ff8405",
          3617 => x"51a5cc3f",
          3618 => x"8285ec08",
          3619 => x"80df3882",
          3620 => x"84d83359",
          3621 => x"78802e89",
          3622 => x"38828490",
          3623 => x"084480cd",
          3624 => x"398284d9",
          3625 => x"33597880",
          3626 => x"2e883882",
          3627 => x"84980844",
          3628 => x"bc398284",
          3629 => x"da335978",
          3630 => x"802e8838",
          3631 => x"8284a008",
          3632 => x"44ab3982",
          3633 => x"84db3359",
          3634 => x"78802e88",
          3635 => x"388284a8",
          3636 => x"08449a39",
          3637 => x"8284d633",
          3638 => x"5978802e",
          3639 => x"88388284",
          3640 => x"b0084489",
          3641 => x"398284c0",
          3642 => x"08fc8005",
          3643 => x"44b43dfe",
          3644 => x"fc1153ff",
          3645 => x"840551a4",
          3646 => x"da3f8285",
          3647 => x"ec0880de",
          3648 => x"388284d8",
          3649 => x"33597880",
          3650 => x"2e893882",
          3651 => x"84940843",
          3652 => x"80cc3982",
          3653 => x"84d93359",
          3654 => x"78802e88",
          3655 => x"3882849c",
          3656 => x"0843bb39",
          3657 => x"8284da33",
          3658 => x"5978802e",
          3659 => x"88388284",
          3660 => x"a40843aa",
          3661 => x"398284db",
          3662 => x"33597880",
          3663 => x"2e883882",
          3664 => x"84ac0843",
          3665 => x"99398284",
          3666 => x"d6335978",
          3667 => x"802e8838",
          3668 => x"8284b408",
          3669 => x"43883982",
          3670 => x"84c00888",
          3671 => x"0543b43d",
          3672 => x"fef81153",
          3673 => x"ff840551",
          3674 => x"a3e93f82",
          3675 => x"85ec0880",
          3676 => x"2ea93880",
          3677 => x"625c5c7a",
          3678 => x"882e8338",
          3679 => x"815c7a90",
          3680 => x"32700981",
          3681 => x"05707207",
          3682 => x"9f2a707f",
          3683 => x"0651515a",
          3684 => x"5a78802e",
          3685 => x"88387aa0",
          3686 => x"2e833888",
          3687 => x"4281f2dc",
          3688 => x"519bc83f",
          3689 => x"a0556354",
          3690 => x"61536252",
          3691 => x"6351f2bf",
          3692 => x"3f81f2ec",
          3693 => x"519bb43f",
          3694 => x"f9d839b4",
          3695 => x"3dff8011",
          3696 => x"53ff8405",
          3697 => x"51a38c3f",
          3698 => x"8285ec08",
          3699 => x"802ef9c2",
          3700 => x"38b43dfe",
          3701 => x"fc1153ff",
          3702 => x"840551a2",
          3703 => x"f63f8285",
          3704 => x"ec08802e",
          3705 => x"a4386359",
          3706 => x"0280cb05",
          3707 => x"33793463",
          3708 => x"810544b4",
          3709 => x"3dfefc11",
          3710 => x"53ff8405",
          3711 => x"51a2d43f",
          3712 => x"8285ec08",
          3713 => x"e138f98a",
          3714 => x"39637033",
          3715 => x"545281f2",
          3716 => x"f851a0c7",
          3717 => x"3f80f852",
          3718 => x"7951a199",
          3719 => x"3f794579",
          3720 => x"335978ae",
          3721 => x"2ef8eb38",
          3722 => x"9f79279f",
          3723 => x"38b43dfe",
          3724 => x"fc1153ff",
          3725 => x"840551a2",
          3726 => x"9a3f8285",
          3727 => x"ec08802e",
          3728 => x"91386359",
          3729 => x"0280cb05",
          3730 => x"33793463",
          3731 => x"810544ff",
          3732 => x"b83981f3",
          3733 => x"84519a93",
          3734 => x"3fffae39",
          3735 => x"b43dfef4",
          3736 => x"1153ff84",
          3737 => x"0551a3e7",
          3738 => x"3f8285ec",
          3739 => x"08802ef8",
          3740 => x"a138b43d",
          3741 => x"fef01153",
          3742 => x"ff840551",
          3743 => x"a3d13f82",
          3744 => x"85ec0880",
          3745 => x"2ea53860",
          3746 => x"5902be05",
          3747 => x"22797082",
          3748 => x"055b2378",
          3749 => x"41b43dfe",
          3750 => x"f01153ff",
          3751 => x"840551a3",
          3752 => x"ae3f8285",
          3753 => x"ec08e038",
          3754 => x"f7e83960",
          3755 => x"70225452",
          3756 => x"81f38c51",
          3757 => x"9fa53f80",
          3758 => x"f8527951",
          3759 => x"9ff73f79",
          3760 => x"45793359",
          3761 => x"78ae2ef7",
          3762 => x"c938789f",
          3763 => x"26873860",
          3764 => x"820541d7",
          3765 => x"39b43dfe",
          3766 => x"f01153ff",
          3767 => x"840551a2",
          3768 => x"ee3f8285",
          3769 => x"ec08802e",
          3770 => x"92386059",
          3771 => x"02be0522",
          3772 => x"79708205",
          3773 => x"5b237841",
          3774 => x"ffb13981",
          3775 => x"f3845198",
          3776 => x"ea3fffa7",
          3777 => x"39b43dfe",
          3778 => x"f41153ff",
          3779 => x"840551a2",
          3780 => x"be3f8285",
          3781 => x"ec08802e",
          3782 => x"f6f838b4",
          3783 => x"3dfef011",
          3784 => x"53ff8405",
          3785 => x"51a2a83f",
          3786 => x"8285ec08",
          3787 => x"802ea038",
          3788 => x"6060710c",
          3789 => x"59608405",
          3790 => x"41b43dfe",
          3791 => x"f01153ff",
          3792 => x"840551a2",
          3793 => x"8a3f8285",
          3794 => x"ec08e538",
          3795 => x"f6c43960",
          3796 => x"70085452",
          3797 => x"81f39851",
          3798 => x"9e813f80",
          3799 => x"f8527951",
          3800 => x"9ed33f79",
          3801 => x"45793359",
          3802 => x"78ae2ef6",
          3803 => x"a5389f79",
          3804 => x"279b38b4",
          3805 => x"3dfef011",
          3806 => x"53ff8405",
          3807 => x"51a1d03f",
          3808 => x"8285ec08",
          3809 => x"802e8d38",
          3810 => x"6060710c",
          3811 => x"59608405",
          3812 => x"41ffbc39",
          3813 => x"81f38451",
          3814 => x"97d13fff",
          3815 => x"b239b43d",
          3816 => x"ff801153",
          3817 => x"ff840551",
          3818 => x"9fa93f82",
          3819 => x"85ec0880",
          3820 => x"2ef5df38",
          3821 => x"635281f3",
          3822 => x"a4519d9f",
          3823 => x"3f635978",
          3824 => x"04b43dff",
          3825 => x"801153ff",
          3826 => x"8405519f",
          3827 => x"863f8285",
          3828 => x"ec08802e",
          3829 => x"f5bc3863",
          3830 => x"5281f3c0",
          3831 => x"519cfc3f",
          3832 => x"6359782d",
          3833 => x"8285ec08",
          3834 => x"802ef5a6",
          3835 => x"388285ec",
          3836 => x"085281f3",
          3837 => x"dc519ce3",
          3838 => x"3ff59739",
          3839 => x"81f3f851",
          3840 => x"96e93fdb",
          3841 => x"963ff58a",
          3842 => x"3981f494",
          3843 => x"5196dc3f",
          3844 => x"8059ffab",
          3845 => x"3990ef3f",
          3846 => x"f4f83979",
          3847 => x"45793359",
          3848 => x"78802ef4",
          3849 => x"ed387d7d",
          3850 => x"06597880",
          3851 => x"2e81d038",
          3852 => x"b43dff84",
          3853 => x"055183b5",
          3854 => x"3f8285ec",
          3855 => x"085c815b",
          3856 => x"7a822eb1",
          3857 => x"387a8224",
          3858 => x"89387a81",
          3859 => x"2e8c3880",
          3860 => x"ca397a83",
          3861 => x"2eae3880",
          3862 => x"c23981f4",
          3863 => x"a8567b55",
          3864 => x"81f4ac54",
          3865 => x"805381f4",
          3866 => x"b052b43d",
          3867 => x"ffb00551",
          3868 => x"9bff3fb8",
          3869 => x"3981f4d0",
          3870 => x"52b43dff",
          3871 => x"b005519b",
          3872 => x"f03fa939",
          3873 => x"7b5581f4",
          3874 => x"ac548053",
          3875 => x"81f4c052",
          3876 => x"b43dffb0",
          3877 => x"05519bd9",
          3878 => x"3f92397b",
          3879 => x"54805381",
          3880 => x"f4cc52b4",
          3881 => x"3dffb005",
          3882 => x"519bc63f",
          3883 => x"82849058",
          3884 => x"8285fc57",
          3885 => x"80566455",
          3886 => x"805482a0",
          3887 => x"805382a0",
          3888 => x"8052b43d",
          3889 => x"ffb00551",
          3890 => x"ebdc3f82",
          3891 => x"85ec0882",
          3892 => x"85ec0809",
          3893 => x"70098105",
          3894 => x"70720780",
          3895 => x"25515b5b",
          3896 => x"5f805a7a",
          3897 => x"83268338",
          3898 => x"815a787a",
          3899 => x"06597880",
          3900 => x"2e8d3881",
          3901 => x"1b7081ff",
          3902 => x"065c597a",
          3903 => x"fec2387d",
          3904 => x"81327d81",
          3905 => x"32075978",
          3906 => x"8a387eff",
          3907 => x"2e098106",
          3908 => x"f3803881",
          3909 => x"f4d4519a",
          3910 => x"c23ff2f6",
          3911 => x"39fc3d0d",
          3912 => x"800b8285",
          3913 => x"fc3487c0",
          3914 => x"948c7008",
          3915 => x"54558784",
          3916 => x"80527251",
          3917 => x"e3d43f82",
          3918 => x"85ec0890",
          3919 => x"2b750855",
          3920 => x"53878480",
          3921 => x"527351e3",
          3922 => x"c13f7282",
          3923 => x"85ec0807",
          3924 => x"750c87c0",
          3925 => x"949c7008",
          3926 => x"54558784",
          3927 => x"80527251",
          3928 => x"e3a83f82",
          3929 => x"85ec0890",
          3930 => x"2b750855",
          3931 => x"53878480",
          3932 => x"527351e3",
          3933 => x"953f7282",
          3934 => x"85ec0807",
          3935 => x"750c8c80",
          3936 => x"830b87c0",
          3937 => x"94840c8c",
          3938 => x"80830b87",
          3939 => x"c094940c",
          3940 => x"80c09a0b",
          3941 => x"829cf40c",
          3942 => x"80c3950b",
          3943 => x"829cf80c",
          3944 => x"89983f92",
          3945 => x"d73f81f4",
          3946 => x"e45193bf",
          3947 => x"3f81f4f0",
          3948 => x"5193b83f",
          3949 => x"a9855192",
          3950 => x"be3f8151",
          3951 => x"ed8c3ff1",
          3952 => x"823f8004",
          3953 => x"fe3d0d80",
          3954 => x"52835371",
          3955 => x"882b5287",
          3956 => x"c43f8285",
          3957 => x"ec0881ff",
          3958 => x"067207ff",
          3959 => x"14545272",
          3960 => x"8025e838",
          3961 => x"718285ec",
          3962 => x"0c843d0d",
          3963 => x"04fc3d0d",
          3964 => x"76700854",
          3965 => x"55807352",
          3966 => x"5472742e",
          3967 => x"818c3872",
          3968 => x"335170a0",
          3969 => x"2e098106",
          3970 => x"86388113",
          3971 => x"53f13972",
          3972 => x"335170a2",
          3973 => x"2e098106",
          3974 => x"86388113",
          3975 => x"53815472",
          3976 => x"5273812e",
          3977 => x"0981069f",
          3978 => x"38843981",
          3979 => x"12528072",
          3980 => x"33525470",
          3981 => x"a22e8338",
          3982 => x"81547080",
          3983 => x"2e9d3873",
          3984 => x"ea389839",
          3985 => x"81125280",
          3986 => x"72335254",
          3987 => x"70a02e83",
          3988 => x"38815470",
          3989 => x"802e8438",
          3990 => x"73ea3880",
          3991 => x"72335254",
          3992 => x"70a02e09",
          3993 => x"81068338",
          3994 => x"815470a2",
          3995 => x"32700981",
          3996 => x"05708025",
          3997 => x"76075151",
          3998 => x"5170802e",
          3999 => x"88388072",
          4000 => x"70810554",
          4001 => x"3471750c",
          4002 => x"72517082",
          4003 => x"85ec0c86",
          4004 => x"3d0d04fc",
          4005 => x"3d0d7653",
          4006 => x"7208802e",
          4007 => x"9138863d",
          4008 => x"fc055272",
          4009 => x"519ba83f",
          4010 => x"8285ec08",
          4011 => x"85388053",
          4012 => x"83397453",
          4013 => x"728285ec",
          4014 => x"0c863d0d",
          4015 => x"04fc3d0d",
          4016 => x"76821133",
          4017 => x"ff055253",
          4018 => x"8152708b",
          4019 => x"26819838",
          4020 => x"831333ff",
          4021 => x"05518252",
          4022 => x"709e2681",
          4023 => x"8a388413",
          4024 => x"33518352",
          4025 => x"70972680",
          4026 => x"fe388513",
          4027 => x"33518452",
          4028 => x"70bb2680",
          4029 => x"f2388613",
          4030 => x"33518552",
          4031 => x"70bb2680",
          4032 => x"e6388813",
          4033 => x"22558652",
          4034 => x"7487e726",
          4035 => x"80d9388a",
          4036 => x"13225487",
          4037 => x"527387e7",
          4038 => x"2680cc38",
          4039 => x"810b87c0",
          4040 => x"989c0c72",
          4041 => x"2287c098",
          4042 => x"bc0c8213",
          4043 => x"3387c098",
          4044 => x"b80c8313",
          4045 => x"3387c098",
          4046 => x"b40c8413",
          4047 => x"3387c098",
          4048 => x"b00c8513",
          4049 => x"3387c098",
          4050 => x"ac0c8613",
          4051 => x"3387c098",
          4052 => x"a80c7487",
          4053 => x"c098a40c",
          4054 => x"7387c098",
          4055 => x"a00c800b",
          4056 => x"87c0989c",
          4057 => x"0c805271",
          4058 => x"8285ec0c",
          4059 => x"863d0d04",
          4060 => x"f33d0d7f",
          4061 => x"5b87c098",
          4062 => x"9c5d817d",
          4063 => x"0c87c098",
          4064 => x"bc085e7d",
          4065 => x"7b2387c0",
          4066 => x"98b8085a",
          4067 => x"79821c34",
          4068 => x"87c098b4",
          4069 => x"085a7983",
          4070 => x"1c3487c0",
          4071 => x"98b0085a",
          4072 => x"79841c34",
          4073 => x"87c098ac",
          4074 => x"085a7985",
          4075 => x"1c3487c0",
          4076 => x"98a8085a",
          4077 => x"79861c34",
          4078 => x"87c098a4",
          4079 => x"085c7b88",
          4080 => x"1c2387c0",
          4081 => x"98a0085a",
          4082 => x"798a1c23",
          4083 => x"807d0c79",
          4084 => x"83ffff06",
          4085 => x"597b83ff",
          4086 => x"ff065886",
          4087 => x"1b335785",
          4088 => x"1b335684",
          4089 => x"1b335583",
          4090 => x"1b335482",
          4091 => x"1b33537d",
          4092 => x"83ffff06",
          4093 => x"5281f588",
          4094 => x"5194e03f",
          4095 => x"8f3d0d04",
          4096 => x"ff3d0d02",
          4097 => x"8f053370",
          4098 => x"09810570",
          4099 => x"9f2a5152",
          4100 => x"52708284",
          4101 => x"8c34833d",
          4102 => x"0d04fb3d",
          4103 => x"0d778284",
          4104 => x"8c337081",
          4105 => x"ff065755",
          4106 => x"5687c094",
          4107 => x"84517480",
          4108 => x"2e863887",
          4109 => x"c0949451",
          4110 => x"70087096",
          4111 => x"2a708106",
          4112 => x"53545270",
          4113 => x"802e8c38",
          4114 => x"71912a70",
          4115 => x"81065151",
          4116 => x"70d73872",
          4117 => x"81327081",
          4118 => x"06515170",
          4119 => x"802e8d38",
          4120 => x"71932a70",
          4121 => x"81065151",
          4122 => x"70ffbe38",
          4123 => x"7381ff06",
          4124 => x"5187c094",
          4125 => x"80527080",
          4126 => x"2e863887",
          4127 => x"c0949052",
          4128 => x"75720c75",
          4129 => x"8285ec0c",
          4130 => x"873d0d04",
          4131 => x"fb3d0d02",
          4132 => x"9f053382",
          4133 => x"848c3370",
          4134 => x"81ff0657",
          4135 => x"555687c0",
          4136 => x"94845174",
          4137 => x"802e8638",
          4138 => x"87c09494",
          4139 => x"51700870",
          4140 => x"962a7081",
          4141 => x"06535452",
          4142 => x"70802e8c",
          4143 => x"3871912a",
          4144 => x"70810651",
          4145 => x"5170d738",
          4146 => x"72813270",
          4147 => x"81065151",
          4148 => x"70802e8d",
          4149 => x"3871932a",
          4150 => x"70810651",
          4151 => x"5170ffbe",
          4152 => x"387381ff",
          4153 => x"065187c0",
          4154 => x"94805270",
          4155 => x"802e8638",
          4156 => x"87c09490",
          4157 => x"5275720c",
          4158 => x"873d0d04",
          4159 => x"f93d0d79",
          4160 => x"54807433",
          4161 => x"7081ff06",
          4162 => x"53535770",
          4163 => x"772e80fc",
          4164 => x"387181ff",
          4165 => x"06811582",
          4166 => x"848c3370",
          4167 => x"81ff0659",
          4168 => x"57555887",
          4169 => x"c0948451",
          4170 => x"75802e86",
          4171 => x"3887c094",
          4172 => x"94517008",
          4173 => x"70962a70",
          4174 => x"81065354",
          4175 => x"5270802e",
          4176 => x"8c387191",
          4177 => x"2a708106",
          4178 => x"515170d7",
          4179 => x"38728132",
          4180 => x"70810651",
          4181 => x"5170802e",
          4182 => x"8d387193",
          4183 => x"2a708106",
          4184 => x"515170ff",
          4185 => x"be387481",
          4186 => x"ff065187",
          4187 => x"c0948052",
          4188 => x"70802e86",
          4189 => x"3887c094",
          4190 => x"90527772",
          4191 => x"0c811774",
          4192 => x"337081ff",
          4193 => x"06535357",
          4194 => x"70ff8638",
          4195 => x"768285ec",
          4196 => x"0c893d0d",
          4197 => x"04fe3d0d",
          4198 => x"82848c33",
          4199 => x"7081ff06",
          4200 => x"545287c0",
          4201 => x"94845172",
          4202 => x"802e8638",
          4203 => x"87c09494",
          4204 => x"51700870",
          4205 => x"822a7081",
          4206 => x"06515151",
          4207 => x"70802ee2",
          4208 => x"387181ff",
          4209 => x"065187c0",
          4210 => x"94805270",
          4211 => x"802e8638",
          4212 => x"87c09490",
          4213 => x"52710870",
          4214 => x"81ff0682",
          4215 => x"85ec0c51",
          4216 => x"843d0d04",
          4217 => x"fe3d0d82",
          4218 => x"848c3370",
          4219 => x"81ff0652",
          4220 => x"5387c094",
          4221 => x"84527080",
          4222 => x"2e863887",
          4223 => x"c0949452",
          4224 => x"71087082",
          4225 => x"2a708106",
          4226 => x"515151ff",
          4227 => x"5270802e",
          4228 => x"a0387281",
          4229 => x"ff065187",
          4230 => x"c0948052",
          4231 => x"70802e86",
          4232 => x"3887c094",
          4233 => x"90527108",
          4234 => x"70982b70",
          4235 => x"982c5153",
          4236 => x"51718285",
          4237 => x"ec0c843d",
          4238 => x"0d04ff3d",
          4239 => x"0d87c09e",
          4240 => x"8008709c",
          4241 => x"2a8a0651",
          4242 => x"5170802e",
          4243 => x"84b43887",
          4244 => x"c09ea408",
          4245 => x"8284900c",
          4246 => x"87c09ea8",
          4247 => x"08828494",
          4248 => x"0c87c09e",
          4249 => x"94088284",
          4250 => x"980c87c0",
          4251 => x"9e980882",
          4252 => x"849c0c87",
          4253 => x"c09e9c08",
          4254 => x"8284a00c",
          4255 => x"87c09ea0",
          4256 => x"088284a4",
          4257 => x"0c87c09e",
          4258 => x"ac088284",
          4259 => x"a80c87c0",
          4260 => x"9eb00882",
          4261 => x"84ac0c87",
          4262 => x"c09eb408",
          4263 => x"8284b00c",
          4264 => x"87c09eb8",
          4265 => x"088284b4",
          4266 => x"0c87c09e",
          4267 => x"bc088284",
          4268 => x"b80c87c0",
          4269 => x"9ec00882",
          4270 => x"84bc0c87",
          4271 => x"c09ec408",
          4272 => x"8284c00c",
          4273 => x"87c09e80",
          4274 => x"08517082",
          4275 => x"84c42387",
          4276 => x"c09e8408",
          4277 => x"8284c80c",
          4278 => x"87c09e88",
          4279 => x"088284cc",
          4280 => x"0c87c09e",
          4281 => x"8c088284",
          4282 => x"d00c810b",
          4283 => x"8284d434",
          4284 => x"800b87c0",
          4285 => x"9e900870",
          4286 => x"84800a06",
          4287 => x"51525270",
          4288 => x"802e8338",
          4289 => x"81527182",
          4290 => x"84d53480",
          4291 => x"0b87c09e",
          4292 => x"90087088",
          4293 => x"800a0651",
          4294 => x"52527080",
          4295 => x"2e833881",
          4296 => x"52718284",
          4297 => x"d634800b",
          4298 => x"87c09e90",
          4299 => x"08709080",
          4300 => x"0a065152",
          4301 => x"5270802e",
          4302 => x"83388152",
          4303 => x"718284d7",
          4304 => x"34800b87",
          4305 => x"c09e9008",
          4306 => x"70888080",
          4307 => x"06515252",
          4308 => x"70802e83",
          4309 => x"38815271",
          4310 => x"8284d834",
          4311 => x"800b87c0",
          4312 => x"9e900870",
          4313 => x"a0808006",
          4314 => x"51525270",
          4315 => x"802e8338",
          4316 => x"81527182",
          4317 => x"84d93480",
          4318 => x"0b87c09e",
          4319 => x"90087090",
          4320 => x"80800651",
          4321 => x"52527080",
          4322 => x"2e833881",
          4323 => x"52718284",
          4324 => x"da34800b",
          4325 => x"87c09e90",
          4326 => x"08708480",
          4327 => x"80065152",
          4328 => x"5270802e",
          4329 => x"83388152",
          4330 => x"718284db",
          4331 => x"34800b87",
          4332 => x"c09e9008",
          4333 => x"70828080",
          4334 => x"06515252",
          4335 => x"70802e83",
          4336 => x"38815271",
          4337 => x"8284dc34",
          4338 => x"800b87c0",
          4339 => x"9e900870",
          4340 => x"81808006",
          4341 => x"51525270",
          4342 => x"802e8338",
          4343 => x"81527182",
          4344 => x"84dd3480",
          4345 => x"0b87c09e",
          4346 => x"90087080",
          4347 => x"c0800651",
          4348 => x"52527080",
          4349 => x"2e833881",
          4350 => x"52718284",
          4351 => x"de34800b",
          4352 => x"87c09e90",
          4353 => x"0870a080",
          4354 => x"06515252",
          4355 => x"70802e83",
          4356 => x"38815271",
          4357 => x"8284df34",
          4358 => x"87c09e90",
          4359 => x"08709880",
          4360 => x"06708a2a",
          4361 => x"51515170",
          4362 => x"8284e034",
          4363 => x"800b87c0",
          4364 => x"9e900870",
          4365 => x"84800651",
          4366 => x"52527080",
          4367 => x"2e833881",
          4368 => x"52718284",
          4369 => x"e13487c0",
          4370 => x"9e900870",
          4371 => x"83f00670",
          4372 => x"842a5151",
          4373 => x"51708284",
          4374 => x"e234800b",
          4375 => x"87c09e90",
          4376 => x"08708806",
          4377 => x"51525270",
          4378 => x"802e8338",
          4379 => x"81527182",
          4380 => x"84e33487",
          4381 => x"c09e9008",
          4382 => x"70870651",
          4383 => x"51708284",
          4384 => x"e434833d",
          4385 => x"0d04fc3d",
          4386 => x"0d81f5a0",
          4387 => x"5185dc3f",
          4388 => x"8284d433",
          4389 => x"5473802e",
          4390 => x"883881f5",
          4391 => x"b45185cb",
          4392 => x"3f81f5c8",
          4393 => x"5185c43f",
          4394 => x"8284d633",
          4395 => x"5473802e",
          4396 => x"93388284",
          4397 => x"b0088284",
          4398 => x"b4081154",
          4399 => x"5281f5e0",
          4400 => x"518b983f",
          4401 => x"8284db33",
          4402 => x"5473802e",
          4403 => x"93388284",
          4404 => x"a8088284",
          4405 => x"ac081154",
          4406 => x"5281f5fc",
          4407 => x"518afc3f",
          4408 => x"8284d833",
          4409 => x"5473802e",
          4410 => x"93388284",
          4411 => x"90088284",
          4412 => x"94081154",
          4413 => x"5281f698",
          4414 => x"518ae03f",
          4415 => x"8284d933",
          4416 => x"5473802e",
          4417 => x"93388284",
          4418 => x"98088284",
          4419 => x"9c081154",
          4420 => x"5281f6b4",
          4421 => x"518ac43f",
          4422 => x"8284da33",
          4423 => x"5473802e",
          4424 => x"93388284",
          4425 => x"a0088284",
          4426 => x"a4081154",
          4427 => x"5281f6d0",
          4428 => x"518aa83f",
          4429 => x"8284df33",
          4430 => x"5473802e",
          4431 => x"8d388284",
          4432 => x"e0335281",
          4433 => x"f6ec518a",
          4434 => x"923f8284",
          4435 => x"e3335473",
          4436 => x"802e8d38",
          4437 => x"8284e433",
          4438 => x"5281f78c",
          4439 => x"5189fc3f",
          4440 => x"8284e133",
          4441 => x"5473802e",
          4442 => x"8d388284",
          4443 => x"e2335281",
          4444 => x"f7ac5189",
          4445 => x"e63f8284",
          4446 => x"d5335473",
          4447 => x"802e8838",
          4448 => x"81f7cc51",
          4449 => x"83e53f82",
          4450 => x"84d73354",
          4451 => x"73802e88",
          4452 => x"3881f7e0",
          4453 => x"5183d43f",
          4454 => x"8284dc33",
          4455 => x"5473802e",
          4456 => x"883881f7",
          4457 => x"ec5183c3",
          4458 => x"3f8284dd",
          4459 => x"33547380",
          4460 => x"2e883881",
          4461 => x"f7f85183",
          4462 => x"b23f8284",
          4463 => x"de335473",
          4464 => x"802e8838",
          4465 => x"81f88451",
          4466 => x"83a13f81",
          4467 => x"f8905183",
          4468 => x"9a3f8284",
          4469 => x"b8085281",
          4470 => x"f89c5188",
          4471 => x"fe3f8284",
          4472 => x"bc085281",
          4473 => x"f8c45188",
          4474 => x"f23f8284",
          4475 => x"c0085281",
          4476 => x"f8ec5188",
          4477 => x"e63f81f9",
          4478 => x"945182ef",
          4479 => x"3f8284c4",
          4480 => x"225281f9",
          4481 => x"9c5188d3",
          4482 => x"3f8284c8",
          4483 => x"0855bd84",
          4484 => x"c0527451",
          4485 => x"d1f43f82",
          4486 => x"85ec0854",
          4487 => x"bd84c052",
          4488 => x"8285ec08",
          4489 => x"51d0e33f",
          4490 => x"748285ec",
          4491 => x"08315373",
          4492 => x"5281f9c4",
          4493 => x"5188a43f",
          4494 => x"8284db33",
          4495 => x"5473802e",
          4496 => x"b0388284",
          4497 => x"cc0855bd",
          4498 => x"84c05274",
          4499 => x"51d1bb3f",
          4500 => x"8285ec08",
          4501 => x"54bd84c0",
          4502 => x"528285ec",
          4503 => x"0851d0aa",
          4504 => x"3f748285",
          4505 => x"ec083153",
          4506 => x"735281f9",
          4507 => x"f05187eb",
          4508 => x"3f8284d6",
          4509 => x"33547380",
          4510 => x"2eb03882",
          4511 => x"84d00855",
          4512 => x"bd84c052",
          4513 => x"7451d182",
          4514 => x"3f8285ec",
          4515 => x"0854bd84",
          4516 => x"c0528285",
          4517 => x"ec0851cf",
          4518 => x"f13f7482",
          4519 => x"85ec0831",
          4520 => x"53735281",
          4521 => x"fa9c5187",
          4522 => x"b23f81f2",
          4523 => x"d85181bb",
          4524 => x"3f863d0d",
          4525 => x"04fe3d0d",
          4526 => x"02920533",
          4527 => x"ff055271",
          4528 => x"8426a938",
          4529 => x"71822b52",
          4530 => x"81e8dc12",
          4531 => x"080481fa",
          4532 => x"c8519d39",
          4533 => x"81fad051",
          4534 => x"973981fa",
          4535 => x"d8519139",
          4536 => x"81fae051",
          4537 => x"8b3981fa",
          4538 => x"e4518539",
          4539 => x"81faec51",
          4540 => x"80f93f84",
          4541 => x"3d0d0471",
          4542 => x"88800c04",
          4543 => x"800b87c0",
          4544 => x"96840c04",
          4545 => x"8284e808",
          4546 => x"87c09684",
          4547 => x"0c04fe3d",
          4548 => x"0d029305",
          4549 => x"3353728a",
          4550 => x"2e098106",
          4551 => x"85388d51",
          4552 => x"ed3f829c",
          4553 => x"fc085271",
          4554 => x"802e9038",
          4555 => x"72723482",
          4556 => x"9cfc0881",
          4557 => x"05829cfc",
          4558 => x"0c8f3982",
          4559 => x"9cf40852",
          4560 => x"71802e85",
          4561 => x"38725171",
          4562 => x"2d843d0d",
          4563 => x"04fe3d0d",
          4564 => x"02970533",
          4565 => x"829cf408",
          4566 => x"76829cf4",
          4567 => x"0c5451ff",
          4568 => x"ad3f7282",
          4569 => x"9cf40c84",
          4570 => x"3d0d04fd",
          4571 => x"3d0d7554",
          4572 => x"73337081",
          4573 => x"ff065353",
          4574 => x"71802e8e",
          4575 => x"387281ff",
          4576 => x"06518114",
          4577 => x"54ff873f",
          4578 => x"e739853d",
          4579 => x"0d04fc3d",
          4580 => x"0d77829c",
          4581 => x"f4087882",
          4582 => x"9cf40c56",
          4583 => x"54733370",
          4584 => x"81ff0653",
          4585 => x"5371802e",
          4586 => x"8e387281",
          4587 => x"ff065181",
          4588 => x"1454feda",
          4589 => x"3fe73974",
          4590 => x"829cf40c",
          4591 => x"863d0d04",
          4592 => x"ec3d0d66",
          4593 => x"68595978",
          4594 => x"7081055a",
          4595 => x"33567580",
          4596 => x"2e858438",
          4597 => x"75a52e09",
          4598 => x"810682e4",
          4599 => x"3880707a",
          4600 => x"7081055c",
          4601 => x"33585b5b",
          4602 => x"75b02e09",
          4603 => x"81068538",
          4604 => x"815a8b39",
          4605 => x"75ad2e09",
          4606 => x"81068a38",
          4607 => x"825a7870",
          4608 => x"81055a33",
          4609 => x"5675aa2e",
          4610 => x"09810692",
          4611 => x"38778419",
          4612 => x"71087b70",
          4613 => x"81055d33",
          4614 => x"595d5953",
          4615 => x"9f39d016",
          4616 => x"53728926",
          4617 => x"97387a83",
          4618 => x"2b7b117c",
          4619 => x"1118d005",
          4620 => x"7b708105",
          4621 => x"5d33595d",
          4622 => x"5153e339",
          4623 => x"7580ec32",
          4624 => x"70098105",
          4625 => x"70720780",
          4626 => x"257880cc",
          4627 => x"32700981",
          4628 => x"05707207",
          4629 => x"80257307",
          4630 => x"53545851",
          4631 => x"55537380",
          4632 => x"2e8c3879",
          4633 => x"84077970",
          4634 => x"81055b33",
          4635 => x"575a7580",
          4636 => x"2e83e438",
          4637 => x"755480e0",
          4638 => x"76278938",
          4639 => x"e0167081",
          4640 => x"ff065553",
          4641 => x"7380cf2e",
          4642 => x"81aa3873",
          4643 => x"80cf24a2",
          4644 => x"387380c3",
          4645 => x"2e818e38",
          4646 => x"7380c324",
          4647 => x"8b387380",
          4648 => x"c22e818c",
          4649 => x"38819939",
          4650 => x"7380c42e",
          4651 => x"818a3881",
          4652 => x"8f397380",
          4653 => x"d52e8180",
          4654 => x"387380d5",
          4655 => x"248a3873",
          4656 => x"80d32e8e",
          4657 => x"3880f939",
          4658 => x"7380d82e",
          4659 => x"80ee3880",
          4660 => x"ef397784",
          4661 => x"19710856",
          4662 => x"59538074",
          4663 => x"33545572",
          4664 => x"752e8d38",
          4665 => x"81157015",
          4666 => x"70335154",
          4667 => x"5572f538",
          4668 => x"79812a56",
          4669 => x"90397481",
          4670 => x"16565372",
          4671 => x"7b278f38",
          4672 => x"a051fc8a",
          4673 => x"3f758106",
          4674 => x"5372802e",
          4675 => x"e9387351",
          4676 => x"fcd93f74",
          4677 => x"81165653",
          4678 => x"727b27fd",
          4679 => x"aa38a051",
          4680 => x"fbec3fef",
          4681 => x"39778419",
          4682 => x"83123353",
          4683 => x"59539339",
          4684 => x"825c9539",
          4685 => x"885c9139",
          4686 => x"8a5c8d39",
          4687 => x"905c8939",
          4688 => x"7551fbca",
          4689 => x"3ffd8039",
          4690 => x"79822a70",
          4691 => x"81065153",
          4692 => x"72802e88",
          4693 => x"38778419",
          4694 => x"59538639",
          4695 => x"84187854",
          4696 => x"58720874",
          4697 => x"80c43270",
          4698 => x"09810570",
          4699 => x"72078025",
          4700 => x"51555555",
          4701 => x"7480258f",
          4702 => x"3872802e",
          4703 => x"8a387409",
          4704 => x"81057a90",
          4705 => x"075b5580",
          4706 => x"0b8f3d5e",
          4707 => x"577b5274",
          4708 => x"51cbaa3f",
          4709 => x"8285ec08",
          4710 => x"81ff067c",
          4711 => x"53755254",
          4712 => x"cae83f82",
          4713 => x"85ec0855",
          4714 => x"89742792",
          4715 => x"38a71453",
          4716 => x"7580f82e",
          4717 => x"84388714",
          4718 => x"537281ff",
          4719 => x"0654b014",
          4720 => x"53727d70",
          4721 => x"81055f34",
          4722 => x"81177509",
          4723 => x"81057077",
          4724 => x"079f2a51",
          4725 => x"5457769f",
          4726 => x"26853872",
          4727 => x"ffaf3879",
          4728 => x"842a7081",
          4729 => x"06515372",
          4730 => x"802e8e38",
          4731 => x"963d7705",
          4732 => x"e00553ad",
          4733 => x"73348117",
          4734 => x"57767a81",
          4735 => x"065455b0",
          4736 => x"54728338",
          4737 => x"a0547981",
          4738 => x"2a708106",
          4739 => x"5456729f",
          4740 => x"38811755",
          4741 => x"767b2797",
          4742 => x"387351f9",
          4743 => x"f13f7581",
          4744 => x"0653728b",
          4745 => x"38748116",
          4746 => x"56537a73",
          4747 => x"26eb3896",
          4748 => x"3d7705e0",
          4749 => x"0553ff17",
          4750 => x"ff147033",
          4751 => x"535457f9",
          4752 => x"cd3f76f2",
          4753 => x"38748116",
          4754 => x"5653727b",
          4755 => x"27faf838",
          4756 => x"a051f9ba",
          4757 => x"3fef3996",
          4758 => x"3d0d04fd",
          4759 => x"3d0d863d",
          4760 => x"70708405",
          4761 => x"52085552",
          4762 => x"7351fad4",
          4763 => x"3f853d0d",
          4764 => x"04fe3d0d",
          4765 => x"74829cfc",
          4766 => x"0c853d88",
          4767 => x"05527551",
          4768 => x"fabe3f82",
          4769 => x"9cfc0853",
          4770 => x"80733480",
          4771 => x"0b829cfc",
          4772 => x"0c843d0d",
          4773 => x"04fd3d0d",
          4774 => x"829cf408",
          4775 => x"76829cf4",
          4776 => x"0c873d88",
          4777 => x"05537752",
          4778 => x"53fa953f",
          4779 => x"72829cf4",
          4780 => x"0c853d0d",
          4781 => x"04fb3d0d",
          4782 => x"7779829c",
          4783 => x"f8087056",
          4784 => x"54575580",
          4785 => x"5471802e",
          4786 => x"80e33882",
          4787 => x"9cf80852",
          4788 => x"712d8285",
          4789 => x"ec0881ff",
          4790 => x"06537280",
          4791 => x"2e80ce38",
          4792 => x"728d2ebc",
          4793 => x"38728832",
          4794 => x"70098105",
          4795 => x"70802551",
          4796 => x"51527380",
          4797 => x"2e8b3871",
          4798 => x"802e8638",
          4799 => x"ff145498",
          4800 => x"399f7325",
          4801 => x"c638ff16",
          4802 => x"52737225",
          4803 => x"ffbd3874",
          4804 => x"14527272",
          4805 => x"34811454",
          4806 => x"7251f7f2",
          4807 => x"3fffac39",
          4808 => x"73155280",
          4809 => x"72348a51",
          4810 => x"f7e43f81",
          4811 => x"53728285",
          4812 => x"ec0c873d",
          4813 => x"0d04fe3d",
          4814 => x"0d829cf8",
          4815 => x"0875829c",
          4816 => x"f80c7753",
          4817 => x"765253fe",
          4818 => x"ec3f7282",
          4819 => x"9cf80c84",
          4820 => x"3d0d04f8",
          4821 => x"3d0d7a7c",
          4822 => x"5a568070",
          4823 => x"7a0c5875",
          4824 => x"08703355",
          4825 => x"5373a02e",
          4826 => x"09810687",
          4827 => x"38811376",
          4828 => x"0ced3973",
          4829 => x"ad2e0981",
          4830 => x"068e3881",
          4831 => x"76081177",
          4832 => x"0c760870",
          4833 => x"33565458",
          4834 => x"73b02e09",
          4835 => x"810680c2",
          4836 => x"38750881",
          4837 => x"05760c75",
          4838 => x"08703355",
          4839 => x"537380e2",
          4840 => x"2e8b3890",
          4841 => x"577380f8",
          4842 => x"2e85388f",
          4843 => x"39825781",
          4844 => x"13760c75",
          4845 => x"08703355",
          4846 => x"53ac3981",
          4847 => x"55a07427",
          4848 => x"818438d0",
          4849 => x"14538055",
          4850 => x"88578973",
          4851 => x"27983880",
          4852 => x"f539d014",
          4853 => x"53805572",
          4854 => x"892680ea",
          4855 => x"38863980",
          4856 => x"5580e339",
          4857 => x"8a578055",
          4858 => x"a0742780",
          4859 => x"ca3880e0",
          4860 => x"74278938",
          4861 => x"e0147081",
          4862 => x"ff065553",
          4863 => x"d0147081",
          4864 => x"ff065553",
          4865 => x"9074278e",
          4866 => x"38f91470",
          4867 => x"81ff0655",
          4868 => x"53897427",
          4869 => x"ca387377",
          4870 => x"27c53876",
          4871 => x"527451c4",
          4872 => x"e93f8285",
          4873 => x"ec081476",
          4874 => x"08810577",
          4875 => x"0c760870",
          4876 => x"33565455",
          4877 => x"ffb23977",
          4878 => x"802e8638",
          4879 => x"74098105",
          4880 => x"5574790c",
          4881 => x"81557482",
          4882 => x"85ec0c8a",
          4883 => x"3d0d04f8",
          4884 => x"3d0d7a7c",
          4885 => x"5a568070",
          4886 => x"7a0c5875",
          4887 => x"08703355",
          4888 => x"5373a02e",
          4889 => x"09810687",
          4890 => x"38811376",
          4891 => x"0ced3973",
          4892 => x"ad2e0981",
          4893 => x"068e3881",
          4894 => x"76081177",
          4895 => x"0c760870",
          4896 => x"33565458",
          4897 => x"73b02e09",
          4898 => x"810680c2",
          4899 => x"38750881",
          4900 => x"05760c75",
          4901 => x"08703355",
          4902 => x"537380e2",
          4903 => x"2e8b3890",
          4904 => x"577380f8",
          4905 => x"2e85388f",
          4906 => x"39825781",
          4907 => x"13760c75",
          4908 => x"08703355",
          4909 => x"53ac3981",
          4910 => x"55a07427",
          4911 => x"818438d0",
          4912 => x"14538055",
          4913 => x"88578973",
          4914 => x"27983880",
          4915 => x"f539d014",
          4916 => x"53805572",
          4917 => x"892680ea",
          4918 => x"38863980",
          4919 => x"5580e339",
          4920 => x"8a578055",
          4921 => x"a0742780",
          4922 => x"ca3880e0",
          4923 => x"74278938",
          4924 => x"e0147081",
          4925 => x"ff065553",
          4926 => x"d0147081",
          4927 => x"ff065553",
          4928 => x"9074278e",
          4929 => x"38f91470",
          4930 => x"81ff0655",
          4931 => x"53897427",
          4932 => x"ca387377",
          4933 => x"27c53876",
          4934 => x"527451c2",
          4935 => x"ed3f8285",
          4936 => x"ec081476",
          4937 => x"08810577",
          4938 => x"0c760870",
          4939 => x"33565455",
          4940 => x"ffb23977",
          4941 => x"802e8638",
          4942 => x"74098105",
          4943 => x"5574790c",
          4944 => x"81557482",
          4945 => x"85ec0c8a",
          4946 => x"3d0d04fd",
          4947 => x"3d0d7698",
          4948 => x"2b70982c",
          4949 => x"79982b70",
          4950 => x"982c7210",
          4951 => x"7311822b",
          4952 => x"54565155",
          4953 => x"5151800b",
          4954 => x"81faf812",
          4955 => x"33555272",
          4956 => x"7425a038",
          4957 => x"7181faf4",
          4958 => x"12081402",
          4959 => x"88059705",
          4960 => x"33713352",
          4961 => x"53535470",
          4962 => x"722e0981",
          4963 => x"06833881",
          4964 => x"54735271",
          4965 => x"8285ec0c",
          4966 => x"853d0d04",
          4967 => x"fc3d0d78",
          4968 => x"0284059f",
          4969 => x"05337133",
          4970 => x"54555371",
          4971 => x"802e9f38",
          4972 => x"8851f2da",
          4973 => x"3fa051f2",
          4974 => x"d53f8851",
          4975 => x"f2d03f72",
          4976 => x"33ff0552",
          4977 => x"71733471",
          4978 => x"81ff0652",
          4979 => x"de397651",
          4980 => x"f3993f73",
          4981 => x"7334863d",
          4982 => x"0d04f63d",
          4983 => x"0d7c0284",
          4984 => x"05b70533",
          4985 => x"028805bb",
          4986 => x"05338285",
          4987 => x"c4337082",
          4988 => x"2b8284ec",
          4989 => x"11085159",
          4990 => x"595a5859",
          4991 => x"74802e86",
          4992 => x"3874519a",
          4993 => x"873f8285",
          4994 => x"c4337082",
          4995 => x"2b8284ec",
          4996 => x"11811a70",
          4997 => x"55595156",
          4998 => x"5a9d883f",
          4999 => x"8285ec08",
          5000 => x"750c8285",
          5001 => x"c4337082",
          5002 => x"2b8284ec",
          5003 => x"11085156",
          5004 => x"5a74802e",
          5005 => x"a7387553",
          5006 => x"78527451",
          5007 => x"ffb8da3f",
          5008 => x"8285c433",
          5009 => x"81055574",
          5010 => x"8285c434",
          5011 => x"7481ff06",
          5012 => x"55937527",
          5013 => x"8738800b",
          5014 => x"8285c434",
          5015 => x"77802eb6",
          5016 => x"388285c0",
          5017 => x"08567580",
          5018 => x"2eac3882",
          5019 => x"85bc3355",
          5020 => x"74a4388c",
          5021 => x"3dfc0554",
          5022 => x"76537852",
          5023 => x"755180d5",
          5024 => x"9f3f8285",
          5025 => x"c008528a",
          5026 => x"51818acd",
          5027 => x"3f8285c0",
          5028 => x"085180d8",
          5029 => x"fc3f8c3d",
          5030 => x"0d04fd3d",
          5031 => x"0d8284ec",
          5032 => x"53935472",
          5033 => x"08527180",
          5034 => x"2e893871",
          5035 => x"5198dd3f",
          5036 => x"80730cff",
          5037 => x"14841454",
          5038 => x"54738025",
          5039 => x"e638800b",
          5040 => x"8285c434",
          5041 => x"8285c008",
          5042 => x"5271802e",
          5043 => x"95387151",
          5044 => x"80d9dc3f",
          5045 => x"8285c008",
          5046 => x"5198b13f",
          5047 => x"800b8285",
          5048 => x"c00c853d",
          5049 => x"0d04dc3d",
          5050 => x"0d815780",
          5051 => x"528285c0",
          5052 => x"085180de",
          5053 => x"c83f8285",
          5054 => x"ec0880d2",
          5055 => x"388285c0",
          5056 => x"085380f8",
          5057 => x"52883d70",
          5058 => x"52568187",
          5059 => x"b33f8285",
          5060 => x"ec08802e",
          5061 => x"b9387551",
          5062 => x"ffb59e3f",
          5063 => x"8285ec08",
          5064 => x"55800b82",
          5065 => x"85ec0825",
          5066 => x"9c388285",
          5067 => x"ec08ff05",
          5068 => x"70175555",
          5069 => x"80743475",
          5070 => x"53765281",
          5071 => x"1781fde8",
          5072 => x"5257f697",
          5073 => x"3f74ff2e",
          5074 => x"098106ff",
          5075 => x"b038a63d",
          5076 => x"0d04d93d",
          5077 => x"0daa3d08",
          5078 => x"ad3d085a",
          5079 => x"5a817058",
          5080 => x"58805282",
          5081 => x"85c00851",
          5082 => x"80ddd23f",
          5083 => x"8285ec08",
          5084 => x"819638ff",
          5085 => x"0b8285c0",
          5086 => x"08545580",
          5087 => x"f8528b3d",
          5088 => x"70525681",
          5089 => x"86ba3f82",
          5090 => x"85ec0880",
          5091 => x"2ea53875",
          5092 => x"51ffb4a5",
          5093 => x"3f8285ec",
          5094 => x"08811858",
          5095 => x"55800b82",
          5096 => x"85ec0825",
          5097 => x"8e388285",
          5098 => x"ec08ff05",
          5099 => x"70175555",
          5100 => x"80743474",
          5101 => x"09700981",
          5102 => x"05707207",
          5103 => x"9f2a5155",
          5104 => x"5578772e",
          5105 => x"853873ff",
          5106 => x"aa388285",
          5107 => x"c0088c11",
          5108 => x"08535180",
          5109 => x"dce73f82",
          5110 => x"85ec0880",
          5111 => x"2e883881",
          5112 => x"fdf451ef",
          5113 => x"863f7877",
          5114 => x"2e098106",
          5115 => x"9b387552",
          5116 => x"7951ffb4",
          5117 => x"b23f7951",
          5118 => x"ffb3be3f",
          5119 => x"ab3d0854",
          5120 => x"8285ec08",
          5121 => x"74348058",
          5122 => x"778285ec",
          5123 => x"0ca93d0d",
          5124 => x"04f63d0d",
          5125 => x"7c7e715c",
          5126 => x"71723357",
          5127 => x"595a5873",
          5128 => x"a02e0981",
          5129 => x"06a23878",
          5130 => x"33780556",
          5131 => x"77762798",
          5132 => x"38811770",
          5133 => x"5b707133",
          5134 => x"56585573",
          5135 => x"a02e0981",
          5136 => x"06863875",
          5137 => x"7526ea38",
          5138 => x"80557483",
          5139 => x"2b8285c8",
          5140 => x"11700853",
          5141 => x"5154ffb2",
          5142 => x"e03f8285",
          5143 => x"ec085379",
          5144 => x"52730851",
          5145 => x"ffb5df3f",
          5146 => x"8285ec08",
          5147 => x"80c33884",
          5148 => x"14335473",
          5149 => x"812e8838",
          5150 => x"73822e88",
          5151 => x"38b339fc",
          5152 => x"e53fbe39",
          5153 => x"811a5a8c",
          5154 => x"3dfc1153",
          5155 => x"f80551f5",
          5156 => x"c23f8285",
          5157 => x"ec08802e",
          5158 => x"9838ff1b",
          5159 => x"53785277",
          5160 => x"51fdaf3f",
          5161 => x"8285ec08",
          5162 => x"81ff0654",
          5163 => x"73802e91",
          5164 => x"38811570",
          5165 => x"81ff0656",
          5166 => x"54827527",
          5167 => x"ff8c3880",
          5168 => x"54738285",
          5169 => x"ec0c8c3d",
          5170 => x"0d04d33d",
          5171 => x"0db03d08",
          5172 => x"b23d08b4",
          5173 => x"3d08595f",
          5174 => x"5a800baf",
          5175 => x"3d348285",
          5176 => x"c4338285",
          5177 => x"c008555b",
          5178 => x"7381ca38",
          5179 => x"738285bc",
          5180 => x"33555573",
          5181 => x"83388155",
          5182 => x"76802e81",
          5183 => x"bb388170",
          5184 => x"76065556",
          5185 => x"73802e81",
          5186 => x"ac38a851",
          5187 => x"97953f82",
          5188 => x"85ec0882",
          5189 => x"85c00c82",
          5190 => x"85ec0880",
          5191 => x"2e819138",
          5192 => x"93537652",
          5193 => x"8285ec08",
          5194 => x"5180c890",
          5195 => x"3f8285ec",
          5196 => x"08802e8b",
          5197 => x"3881fea0",
          5198 => x"51f2a03f",
          5199 => x"80f73982",
          5200 => x"85ec085b",
          5201 => x"8285c008",
          5202 => x"5380f852",
          5203 => x"903d7052",
          5204 => x"548182ec",
          5205 => x"3f8285ec",
          5206 => x"08568285",
          5207 => x"ec08742e",
          5208 => x"09810680",
          5209 => x"d0388285",
          5210 => x"ec0851ff",
          5211 => x"b0cb3f82",
          5212 => x"85ec0855",
          5213 => x"800b8285",
          5214 => x"ec0825a9",
          5215 => x"388285ec",
          5216 => x"08ff0570",
          5217 => x"17555580",
          5218 => x"74348053",
          5219 => x"7481ff06",
          5220 => x"527551f8",
          5221 => x"c53f811b",
          5222 => x"7081ff06",
          5223 => x"5c54937b",
          5224 => x"27833880",
          5225 => x"5b74ff2e",
          5226 => x"098106ff",
          5227 => x"97388639",
          5228 => x"758285bc",
          5229 => x"34768c38",
          5230 => x"8285c008",
          5231 => x"802e8438",
          5232 => x"f9d83f8f",
          5233 => x"3d5de09c",
          5234 => x"3f8285ec",
          5235 => x"08982b70",
          5236 => x"982c5159",
          5237 => x"78ff2eee",
          5238 => x"387881ff",
          5239 => x"06829d84",
          5240 => x"3370982b",
          5241 => x"70982c82",
          5242 => x"9d803370",
          5243 => x"982b7097",
          5244 => x"2c71982c",
          5245 => x"0570822b",
          5246 => x"81faf411",
          5247 => x"08157033",
          5248 => x"51515151",
          5249 => x"59595159",
          5250 => x"5d588156",
          5251 => x"73782e80",
          5252 => x"e3387774",
          5253 => x"27b138ff",
          5254 => x"1570982b",
          5255 => x"70982c51",
          5256 => x"56548075",
          5257 => x"2480cb38",
          5258 => x"76537452",
          5259 => x"7751f69b",
          5260 => x"3f8285ec",
          5261 => x"0881ff06",
          5262 => x"5473802e",
          5263 => x"da387482",
          5264 => x"9d803481",
          5265 => x"56ae3981",
          5266 => x"1570982b",
          5267 => x"70982c70",
          5268 => x"81ff0653",
          5269 => x"51565473",
          5270 => x"95269738",
          5271 => x"76537452",
          5272 => x"7751f5e7",
          5273 => x"3f8285ec",
          5274 => x"0881ff06",
          5275 => x"5473cf38",
          5276 => x"d6398056",
          5277 => x"75802e80",
          5278 => x"ca38811c",
          5279 => x"5473829d",
          5280 => x"84347398",
          5281 => x"2b70982c",
          5282 => x"829d8033",
          5283 => x"70982b70",
          5284 => x"982c7010",
          5285 => x"7111822b",
          5286 => x"81faf811",
          5287 => x"335e5253",
          5288 => x"51585851",
          5289 => x"5473772e",
          5290 => x"098106fe",
          5291 => x"993881fa",
          5292 => x"fc15087d",
          5293 => x"0c800b82",
          5294 => x"9d843480",
          5295 => x"0b829d80",
          5296 => x"34923975",
          5297 => x"829d8434",
          5298 => x"75829d80",
          5299 => x"3478af3d",
          5300 => x"34757d0c",
          5301 => x"7e547395",
          5302 => x"26fde838",
          5303 => x"73822b54",
          5304 => x"81e8f014",
          5305 => x"0804829d",
          5306 => x"8c335675",
          5307 => x"7e2efdd3",
          5308 => x"38829d88",
          5309 => x"33547574",
          5310 => x"27ab3873",
          5311 => x"982b7098",
          5312 => x"2c515575",
          5313 => x"75249e38",
          5314 => x"741a5473",
          5315 => x"33811534",
          5316 => x"ff157098",
          5317 => x"2b70982c",
          5318 => x"829d8c33",
          5319 => x"53515654",
          5320 => x"747425e4",
          5321 => x"38829d8c",
          5322 => x"33811156",
          5323 => x"5474829d",
          5324 => x"8c34731a",
          5325 => x"54ae3d33",
          5326 => x"7434829d",
          5327 => x"88335473",
          5328 => x"7e258938",
          5329 => x"81145473",
          5330 => x"829d8834",
          5331 => x"829d8c33",
          5332 => x"ff057098",
          5333 => x"2b70982c",
          5334 => x"829d8833",
          5335 => x"59515654",
          5336 => x"7476259f",
          5337 => x"38741a70",
          5338 => x"335254e7",
          5339 => x"a13f8115",
          5340 => x"70982b70",
          5341 => x"982c829d",
          5342 => x"88335a51",
          5343 => x"56547675",
          5344 => x"24e33882",
          5345 => x"9d8c3370",
          5346 => x"982b7098",
          5347 => x"2c829d88",
          5348 => x"33595156",
          5349 => x"54747625",
          5350 => x"fca93888",
          5351 => x"51e6ef3f",
          5352 => x"81157098",
          5353 => x"2b70982c",
          5354 => x"829d8833",
          5355 => x"5a515654",
          5356 => x"767524e7",
          5357 => x"38fc8c39",
          5358 => x"837a3480",
          5359 => x"0b811b34",
          5360 => x"829d8c53",
          5361 => x"805281f3",
          5362 => x"d851f3d0",
          5363 => x"3f81d939",
          5364 => x"829d8c33",
          5365 => x"7081ff06",
          5366 => x"55557380",
          5367 => x"2efbe438",
          5368 => x"829d8833",
          5369 => x"ff055473",
          5370 => x"829d8834",
          5371 => x"ff155473",
          5372 => x"829d8c34",
          5373 => x"8851e696",
          5374 => x"3f829d8c",
          5375 => x"3370982b",
          5376 => x"70982c82",
          5377 => x"9d883357",
          5378 => x"51565774",
          5379 => x"7425a438",
          5380 => x"741a5481",
          5381 => x"14337434",
          5382 => x"733351e5",
          5383 => x"f13f8115",
          5384 => x"70982b70",
          5385 => x"982c829d",
          5386 => x"88335951",
          5387 => x"56547575",
          5388 => x"24de38a0",
          5389 => x"51e5d73f",
          5390 => x"829d8c33",
          5391 => x"70982b70",
          5392 => x"982c829d",
          5393 => x"88335751",
          5394 => x"56577474",
          5395 => x"24faf438",
          5396 => x"8851e5ba",
          5397 => x"3f811570",
          5398 => x"982b7098",
          5399 => x"2c829d88",
          5400 => x"33595156",
          5401 => x"54757525",
          5402 => x"e738fad7",
          5403 => x"39829d88",
          5404 => x"337a0554",
          5405 => x"8074348a",
          5406 => x"51e5933f",
          5407 => x"829d8852",
          5408 => x"7951f78d",
          5409 => x"3f8285ec",
          5410 => x"0881ff06",
          5411 => x"54739638",
          5412 => x"829d8833",
          5413 => x"5473802e",
          5414 => x"8f388153",
          5415 => x"73527951",
          5416 => x"f2b83f84",
          5417 => x"39807a34",
          5418 => x"800b829d",
          5419 => x"8c34800b",
          5420 => x"829d8834",
          5421 => x"798285ec",
          5422 => x"0caf3d0d",
          5423 => x"04829d8c",
          5424 => x"33547380",
          5425 => x"2ef9fc38",
          5426 => x"8851e4c2",
          5427 => x"3f829d8c",
          5428 => x"33ff0554",
          5429 => x"73829d8c",
          5430 => x"347381ff",
          5431 => x"0654e339",
          5432 => x"829d8c33",
          5433 => x"829d8833",
          5434 => x"55557375",
          5435 => x"2ef9d438",
          5436 => x"ff145473",
          5437 => x"829d8834",
          5438 => x"74982b70",
          5439 => x"982c7581",
          5440 => x"ff065651",
          5441 => x"55747425",
          5442 => x"a438741a",
          5443 => x"54811433",
          5444 => x"74347333",
          5445 => x"51e3f73f",
          5446 => x"81157098",
          5447 => x"2b70982c",
          5448 => x"829d8833",
          5449 => x"59515654",
          5450 => x"757524de",
          5451 => x"38a051e3",
          5452 => x"dd3f829d",
          5453 => x"8c337098",
          5454 => x"2b70982c",
          5455 => x"829d8833",
          5456 => x"57515657",
          5457 => x"747424f8",
          5458 => x"fa388851",
          5459 => x"e3c03f81",
          5460 => x"1570982b",
          5461 => x"70982c82",
          5462 => x"9d883359",
          5463 => x"51565475",
          5464 => x"7525e738",
          5465 => x"f8dd3982",
          5466 => x"9d8c3370",
          5467 => x"81ff0682",
          5468 => x"9d883359",
          5469 => x"56547477",
          5470 => x"27f8c838",
          5471 => x"81145473",
          5472 => x"829d8c34",
          5473 => x"741a7033",
          5474 => x"5254e382",
          5475 => x"3f829d8c",
          5476 => x"337081ff",
          5477 => x"06829d88",
          5478 => x"33585654",
          5479 => x"757526dc",
          5480 => x"38f8a039",
          5481 => x"829d8c53",
          5482 => x"805281f3",
          5483 => x"d851efec",
          5484 => x"3f800b82",
          5485 => x"9d8c3480",
          5486 => x"0b829d88",
          5487 => x"34f88439",
          5488 => x"7ab03882",
          5489 => x"85b80855",
          5490 => x"74802ea6",
          5491 => x"387451ff",
          5492 => x"a7e73f82",
          5493 => x"85ec0882",
          5494 => x"9d883482",
          5495 => x"85ec0881",
          5496 => x"ff068105",
          5497 => x"53745279",
          5498 => x"51ffa9ad",
          5499 => x"3f935b81",
          5500 => x"c0397a82",
          5501 => x"2b8284ec",
          5502 => x"11fc1108",
          5503 => x"57515474",
          5504 => x"802ea738",
          5505 => x"7451ffa7",
          5506 => x"b03f8285",
          5507 => x"ec08829d",
          5508 => x"88348285",
          5509 => x"ec0881ff",
          5510 => x"06810553",
          5511 => x"74527951",
          5512 => x"ffa8f63f",
          5513 => x"ff1b5480",
          5514 => x"f9397308",
          5515 => x"5574802e",
          5516 => x"f7913874",
          5517 => x"51ffa781",
          5518 => x"3f99397a",
          5519 => x"932e0981",
          5520 => x"06ae3882",
          5521 => x"84ec0855",
          5522 => x"74802ea4",
          5523 => x"387451ff",
          5524 => x"a6e73f82",
          5525 => x"85ec0882",
          5526 => x"9d883482",
          5527 => x"85ec0881",
          5528 => x"ff068105",
          5529 => x"53745279",
          5530 => x"51ffa8ad",
          5531 => x"3f80c239",
          5532 => x"7a822b82",
          5533 => x"84f01108",
          5534 => x"56547480",
          5535 => x"2eab3874",
          5536 => x"51ffa6b5",
          5537 => x"3f8285ec",
          5538 => x"08829d88",
          5539 => x"348285ec",
          5540 => x"0881ff06",
          5541 => x"81055374",
          5542 => x"527951ff",
          5543 => x"a7fb3f81",
          5544 => x"1b547381",
          5545 => x"ff065b89",
          5546 => x"3974829d",
          5547 => x"8834747a",
          5548 => x"34829d8c",
          5549 => x"53829d88",
          5550 => x"33527951",
          5551 => x"edde3ff6",
          5552 => x"8239829d",
          5553 => x"8c337081",
          5554 => x"ff06829d",
          5555 => x"88335956",
          5556 => x"54747727",
          5557 => x"f5ed3881",
          5558 => x"14547382",
          5559 => x"9d8c3474",
          5560 => x"1a703352",
          5561 => x"54e0a73f",
          5562 => x"f5d93982",
          5563 => x"9d8c3354",
          5564 => x"73802ef5",
          5565 => x"ce388851",
          5566 => x"e0943f82",
          5567 => x"9d8c33ff",
          5568 => x"05547382",
          5569 => x"9d8c34f5",
          5570 => x"ba39f93d",
          5571 => x"0d83dff4",
          5572 => x"0b8285e4",
          5573 => x"0c82800b",
          5574 => x"8285e023",
          5575 => x"90805380",
          5576 => x"5283dff4",
          5577 => x"51ffaac5",
          5578 => x"3f8285e4",
          5579 => x"08548058",
          5580 => x"77743481",
          5581 => x"57768115",
          5582 => x"348285e4",
          5583 => x"08547784",
          5584 => x"15347685",
          5585 => x"15348285",
          5586 => x"e4085477",
          5587 => x"86153476",
          5588 => x"87153482",
          5589 => x"85e40882",
          5590 => x"85e022ff",
          5591 => x"05fe8080",
          5592 => x"077083ff",
          5593 => x"ff067088",
          5594 => x"2a585155",
          5595 => x"56748817",
          5596 => x"34738917",
          5597 => x"348285e0",
          5598 => x"2270832b",
          5599 => x"8285e408",
          5600 => x"11f80551",
          5601 => x"55557782",
          5602 => x"15347683",
          5603 => x"1534893d",
          5604 => x"0d04ff3d",
          5605 => x"0d735281",
          5606 => x"51847227",
          5607 => x"8f38fb12",
          5608 => x"832a8211",
          5609 => x"7083ffff",
          5610 => x"06515151",
          5611 => x"708285ec",
          5612 => x"0c833d0d",
          5613 => x"04f93d0d",
          5614 => x"02a60522",
          5615 => x"028405aa",
          5616 => x"05227105",
          5617 => x"8285e408",
          5618 => x"71832b71",
          5619 => x"1174832b",
          5620 => x"73117033",
          5621 => x"81123371",
          5622 => x"882b0702",
          5623 => x"a405ae05",
          5624 => x"227181ff",
          5625 => x"ff060770",
          5626 => x"882a5351",
          5627 => x"5259545b",
          5628 => x"5b575354",
          5629 => x"55717734",
          5630 => x"70811834",
          5631 => x"8285e408",
          5632 => x"1475882a",
          5633 => x"52547082",
          5634 => x"15347483",
          5635 => x"15348285",
          5636 => x"e4087017",
          5637 => x"70338112",
          5638 => x"3371882b",
          5639 => x"0770832b",
          5640 => x"8ffff806",
          5641 => x"51525652",
          5642 => x"71057383",
          5643 => x"ffff0670",
          5644 => x"882a5454",
          5645 => x"51718212",
          5646 => x"347281ff",
          5647 => x"06537283",
          5648 => x"12348285",
          5649 => x"e4081656",
          5650 => x"71763472",
          5651 => x"81173489",
          5652 => x"3d0d04fb",
          5653 => x"3d0d8285",
          5654 => x"e4080284",
          5655 => x"059e0522",
          5656 => x"70832b72",
          5657 => x"11861133",
          5658 => x"87123371",
          5659 => x"8b2b7183",
          5660 => x"2b07585b",
          5661 => x"59525552",
          5662 => x"72058412",
          5663 => x"33851333",
          5664 => x"71882b07",
          5665 => x"70882a54",
          5666 => x"56565270",
          5667 => x"84133473",
          5668 => x"85133482",
          5669 => x"85e40870",
          5670 => x"14841133",
          5671 => x"85123371",
          5672 => x"8b2b7183",
          5673 => x"2b075659",
          5674 => x"57527205",
          5675 => x"86123387",
          5676 => x"13337188",
          5677 => x"2b077088",
          5678 => x"2a545656",
          5679 => x"52708613",
          5680 => x"34738713",
          5681 => x"348285e4",
          5682 => x"08137033",
          5683 => x"81123371",
          5684 => x"882b0770",
          5685 => x"81ffff06",
          5686 => x"70882a53",
          5687 => x"51535353",
          5688 => x"71733470",
          5689 => x"81143487",
          5690 => x"3d0d04f9",
          5691 => x"3d0d02a6",
          5692 => x"05228285",
          5693 => x"e4087183",
          5694 => x"2b711170",
          5695 => x"33811233",
          5696 => x"71882b07",
          5697 => x"70832b53",
          5698 => x"595b5558",
          5699 => x"73057033",
          5700 => x"81123371",
          5701 => x"982b7190",
          5702 => x"2b07535a",
          5703 => x"55535571",
          5704 => x"802580f6",
          5705 => x"387351fe",
          5706 => x"aa3f8285",
          5707 => x"e4087017",
          5708 => x"70338112",
          5709 => x"33718b2b",
          5710 => x"71832b07",
          5711 => x"74117033",
          5712 => x"81123371",
          5713 => x"882b0770",
          5714 => x"832b8fff",
          5715 => x"f8065152",
          5716 => x"5d515357",
          5717 => x"5a537205",
          5718 => x"75882a54",
          5719 => x"52728213",
          5720 => x"34748313",
          5721 => x"348285e4",
          5722 => x"08701770",
          5723 => x"33811233",
          5724 => x"718b2b71",
          5725 => x"832b0756",
          5726 => x"59575572",
          5727 => x"05703381",
          5728 => x"12337188",
          5729 => x"2b077081",
          5730 => x"ffff0670",
          5731 => x"882a5751",
          5732 => x"52585272",
          5733 => x"74347181",
          5734 => x"1534893d",
          5735 => x"0d04fb3d",
          5736 => x"0d8285e4",
          5737 => x"08028405",
          5738 => x"9e052270",
          5739 => x"832b7211",
          5740 => x"82113383",
          5741 => x"1233718b",
          5742 => x"2b71832b",
          5743 => x"07595b59",
          5744 => x"52565273",
          5745 => x"05713381",
          5746 => x"13337188",
          5747 => x"2b07028c",
          5748 => x"05a20522",
          5749 => x"71077088",
          5750 => x"2a535153",
          5751 => x"53537173",
          5752 => x"34708114",
          5753 => x"348285e4",
          5754 => x"08701570",
          5755 => x"33811233",
          5756 => x"718b2b71",
          5757 => x"832b0756",
          5758 => x"59575272",
          5759 => x"05821233",
          5760 => x"83133371",
          5761 => x"882b0770",
          5762 => x"882a5455",
          5763 => x"56527082",
          5764 => x"13347283",
          5765 => x"13348285",
          5766 => x"e4081482",
          5767 => x"11338312",
          5768 => x"3371882b",
          5769 => x"078285ec",
          5770 => x"0c525487",
          5771 => x"3d0d04f7",
          5772 => x"3d0d7b82",
          5773 => x"85e40831",
          5774 => x"832a7083",
          5775 => x"ffff0670",
          5776 => x"535753fd",
          5777 => x"a63f8285",
          5778 => x"e4087683",
          5779 => x"2b711182",
          5780 => x"11338312",
          5781 => x"33718b2b",
          5782 => x"71832b07",
          5783 => x"75117033",
          5784 => x"81123371",
          5785 => x"982b7190",
          5786 => x"2b075342",
          5787 => x"4051535b",
          5788 => x"58555954",
          5789 => x"7280258d",
          5790 => x"38828080",
          5791 => x"527551fe",
          5792 => x"9d3f8184",
          5793 => x"39841433",
          5794 => x"85153371",
          5795 => x"8b2b7183",
          5796 => x"2b077611",
          5797 => x"79882a53",
          5798 => x"51555855",
          5799 => x"76861434",
          5800 => x"7581ff06",
          5801 => x"56758714",
          5802 => x"348285e4",
          5803 => x"08701984",
          5804 => x"12338513",
          5805 => x"3371882b",
          5806 => x"0770882a",
          5807 => x"54575b56",
          5808 => x"53728416",
          5809 => x"34738516",
          5810 => x"348285e4",
          5811 => x"08185380",
          5812 => x"0b861434",
          5813 => x"800b8714",
          5814 => x"348285e4",
          5815 => x"08537684",
          5816 => x"14347585",
          5817 => x"14348285",
          5818 => x"e4081870",
          5819 => x"33811233",
          5820 => x"71882b07",
          5821 => x"70828080",
          5822 => x"0770882a",
          5823 => x"53515556",
          5824 => x"54747434",
          5825 => x"72811534",
          5826 => x"8b3d0d04",
          5827 => x"ff3d0d73",
          5828 => x"528285e4",
          5829 => x"088438f7",
          5830 => x"f13f7180",
          5831 => x"2e863871",
          5832 => x"51fe8c3f",
          5833 => x"833d0d04",
          5834 => x"f53d0d80",
          5835 => x"7e5258f8",
          5836 => x"e13f8285",
          5837 => x"ec0883ff",
          5838 => x"ff068285",
          5839 => x"e4088411",
          5840 => x"33851233",
          5841 => x"71882b07",
          5842 => x"705f5956",
          5843 => x"585a81ff",
          5844 => x"ff597578",
          5845 => x"2e80cc38",
          5846 => x"75832b77",
          5847 => x"05703381",
          5848 => x"12337188",
          5849 => x"2b077081",
          5850 => x"ffff0679",
          5851 => x"317083ff",
          5852 => x"ff06707f",
          5853 => x"27525351",
          5854 => x"56595577",
          5855 => x"79278a38",
          5856 => x"73802e85",
          5857 => x"3875785a",
          5858 => x"5b841533",
          5859 => x"85163371",
          5860 => x"882b0757",
          5861 => x"5475c138",
          5862 => x"7881ffff",
          5863 => x"2e85387a",
          5864 => x"79595680",
          5865 => x"76832b82",
          5866 => x"85e40811",
          5867 => x"70338112",
          5868 => x"3371882b",
          5869 => x"077081ff",
          5870 => x"ff065152",
          5871 => x"5a565c55",
          5872 => x"73752e83",
          5873 => x"38815580",
          5874 => x"54797826",
          5875 => x"81cc3874",
          5876 => x"5474802e",
          5877 => x"81c43877",
          5878 => x"7a2e0981",
          5879 => x"06893875",
          5880 => x"51f8f03f",
          5881 => x"81ac3982",
          5882 => x"80805379",
          5883 => x"527551f7",
          5884 => x"c43f8285",
          5885 => x"e408701c",
          5886 => x"86113387",
          5887 => x"1233718b",
          5888 => x"2b71832b",
          5889 => x"07535a5e",
          5890 => x"5574057a",
          5891 => x"177083ff",
          5892 => x"ff067088",
          5893 => x"2a5c5956",
          5894 => x"54788415",
          5895 => x"347681ff",
          5896 => x"06577685",
          5897 => x"15348285",
          5898 => x"e4087583",
          5899 => x"2b711172",
          5900 => x"1e861133",
          5901 => x"87123371",
          5902 => x"882b0770",
          5903 => x"882a535b",
          5904 => x"5e535a56",
          5905 => x"54738619",
          5906 => x"34758719",
          5907 => x"348285e4",
          5908 => x"08701c84",
          5909 => x"11338512",
          5910 => x"33718b2b",
          5911 => x"71832b07",
          5912 => x"535d5a55",
          5913 => x"74055478",
          5914 => x"86153476",
          5915 => x"87153482",
          5916 => x"85e40870",
          5917 => x"16711d84",
          5918 => x"11338512",
          5919 => x"3371882b",
          5920 => x"0770882a",
          5921 => x"535a5f52",
          5922 => x"56547384",
          5923 => x"16347585",
          5924 => x"16348285",
          5925 => x"e4081b84",
          5926 => x"05547382",
          5927 => x"85ec0c8d",
          5928 => x"3d0d04fe",
          5929 => x"3d0d7452",
          5930 => x"8285e408",
          5931 => x"8438f4da",
          5932 => x"3f715371",
          5933 => x"802e8b38",
          5934 => x"7151fcec",
          5935 => x"3f8285ec",
          5936 => x"08537282",
          5937 => x"85ec0c84",
          5938 => x"3d0d04ff",
          5939 => x"3d0d028f",
          5940 => x"05335181",
          5941 => x"52707226",
          5942 => x"87388285",
          5943 => x"e8113352",
          5944 => x"718285ec",
          5945 => x"0c833d0d",
          5946 => x"04fc3d0d",
          5947 => x"029b0533",
          5948 => x"0284059f",
          5949 => x"05335653",
          5950 => x"83517281",
          5951 => x"2680e038",
          5952 => x"72842b87",
          5953 => x"c0928c11",
          5954 => x"53518854",
          5955 => x"74802e84",
          5956 => x"38818854",
          5957 => x"73720c87",
          5958 => x"c0928c11",
          5959 => x"5181710c",
          5960 => x"850b87c0",
          5961 => x"988c0c70",
          5962 => x"52710870",
          5963 => x"82065151",
          5964 => x"70802e8a",
          5965 => x"3887c098",
          5966 => x"8c085170",
          5967 => x"ec387108",
          5968 => x"fc808006",
          5969 => x"52719238",
          5970 => x"87c0988c",
          5971 => x"08517080",
          5972 => x"2e873871",
          5973 => x"8285e814",
          5974 => x"348285e8",
          5975 => x"13335170",
          5976 => x"8285ec0c",
          5977 => x"863d0d04",
          5978 => x"f33d0d60",
          5979 => x"6264028c",
          5980 => x"05bf0533",
          5981 => x"5740585b",
          5982 => x"8374525a",
          5983 => x"fecd3f82",
          5984 => x"85ec0881",
          5985 => x"067a5452",
          5986 => x"7181be38",
          5987 => x"71727584",
          5988 => x"2b87c092",
          5989 => x"801187c0",
          5990 => x"928c1287",
          5991 => x"c0928413",
          5992 => x"415a4057",
          5993 => x"5a58850b",
          5994 => x"87c0988c",
          5995 => x"0c767d0c",
          5996 => x"84760c75",
          5997 => x"0870852a",
          5998 => x"70810651",
          5999 => x"53547180",
          6000 => x"2e8e387b",
          6001 => x"0852717b",
          6002 => x"7081055d",
          6003 => x"34811959",
          6004 => x"8074a206",
          6005 => x"53537173",
          6006 => x"2e833881",
          6007 => x"537883ff",
          6008 => x"268f3872",
          6009 => x"802e8a38",
          6010 => x"87c0988c",
          6011 => x"085271c3",
          6012 => x"3887c098",
          6013 => x"8c085271",
          6014 => x"802e8738",
          6015 => x"7884802e",
          6016 => x"99388176",
          6017 => x"0c87c092",
          6018 => x"8c155372",
          6019 => x"08708206",
          6020 => x"515271f7",
          6021 => x"38ff1a5a",
          6022 => x"8d398480",
          6023 => x"17811970",
          6024 => x"81ff065a",
          6025 => x"53577980",
          6026 => x"2e903873",
          6027 => x"fc808006",
          6028 => x"52718738",
          6029 => x"7d7826fe",
          6030 => x"ed3873fc",
          6031 => x"80800652",
          6032 => x"71802e83",
          6033 => x"38815271",
          6034 => x"53728285",
          6035 => x"ec0c8f3d",
          6036 => x"0d04f33d",
          6037 => x"0d606264",
          6038 => x"028c05bf",
          6039 => x"05335740",
          6040 => x"585b8359",
          6041 => x"80745258",
          6042 => x"fce13f82",
          6043 => x"85ec0881",
          6044 => x"06795452",
          6045 => x"71782e09",
          6046 => x"810681b1",
          6047 => x"38777484",
          6048 => x"2b87c092",
          6049 => x"801187c0",
          6050 => x"928c1287",
          6051 => x"c0928413",
          6052 => x"40595f56",
          6053 => x"5a850b87",
          6054 => x"c0988c0c",
          6055 => x"767d0c82",
          6056 => x"760c8058",
          6057 => x"75087084",
          6058 => x"2a708106",
          6059 => x"51535471",
          6060 => x"802e8c38",
          6061 => x"7a708105",
          6062 => x"5c337c0c",
          6063 => x"81185873",
          6064 => x"812a7081",
          6065 => x"06515271",
          6066 => x"802e8a38",
          6067 => x"87c0988c",
          6068 => x"085271d0",
          6069 => x"3887c098",
          6070 => x"8c085271",
          6071 => x"802e8738",
          6072 => x"7784802e",
          6073 => x"99388176",
          6074 => x"0c87c092",
          6075 => x"8c155372",
          6076 => x"08708206",
          6077 => x"515271f7",
          6078 => x"38ff1959",
          6079 => x"8d39811a",
          6080 => x"7081ff06",
          6081 => x"84801959",
          6082 => x"5b527880",
          6083 => x"2e903873",
          6084 => x"fc808006",
          6085 => x"52718738",
          6086 => x"7d7a26fe",
          6087 => x"f83873fc",
          6088 => x"80800652",
          6089 => x"71802e83",
          6090 => x"38815271",
          6091 => x"53728285",
          6092 => x"ec0c8f3d",
          6093 => x"0d04fa3d",
          6094 => x"0d7a0284",
          6095 => x"05a30533",
          6096 => x"028805a7",
          6097 => x"05337154",
          6098 => x"545657fa",
          6099 => x"fe3f8285",
          6100 => x"ec088106",
          6101 => x"53835472",
          6102 => x"80fe3885",
          6103 => x"0b87c098",
          6104 => x"8c0c8156",
          6105 => x"71762e80",
          6106 => x"dc387176",
          6107 => x"24933874",
          6108 => x"842b87c0",
          6109 => x"928c1154",
          6110 => x"5471802e",
          6111 => x"8d3880d4",
          6112 => x"3971832e",
          6113 => x"80c63880",
          6114 => x"cb397208",
          6115 => x"70812a70",
          6116 => x"81065151",
          6117 => x"5271802e",
          6118 => x"8a3887c0",
          6119 => x"988c0852",
          6120 => x"71e83887",
          6121 => x"c0988c08",
          6122 => x"52719638",
          6123 => x"81730c87",
          6124 => x"c0928c14",
          6125 => x"53720870",
          6126 => x"82065152",
          6127 => x"71f73896",
          6128 => x"39805692",
          6129 => x"3988800a",
          6130 => x"770c8539",
          6131 => x"8180770c",
          6132 => x"72568339",
          6133 => x"84567554",
          6134 => x"738285ec",
          6135 => x"0c883d0d",
          6136 => x"04fe3d0d",
          6137 => x"74811133",
          6138 => x"71337188",
          6139 => x"2b078285",
          6140 => x"ec0c5351",
          6141 => x"843d0d04",
          6142 => x"fd3d0d75",
          6143 => x"83113382",
          6144 => x"12337190",
          6145 => x"2b71882b",
          6146 => x"07811433",
          6147 => x"70720788",
          6148 => x"2b753371",
          6149 => x"078285ec",
          6150 => x"0c525354",
          6151 => x"56545285",
          6152 => x"3d0d04ff",
          6153 => x"3d0d7302",
          6154 => x"84059205",
          6155 => x"22525270",
          6156 => x"72708105",
          6157 => x"54347088",
          6158 => x"2a517072",
          6159 => x"34833d0d",
          6160 => x"04ff3d0d",
          6161 => x"73755252",
          6162 => x"70727081",
          6163 => x"05543470",
          6164 => x"882a5170",
          6165 => x"72708105",
          6166 => x"54347088",
          6167 => x"2a517072",
          6168 => x"70810554",
          6169 => x"3470882a",
          6170 => x"51707234",
          6171 => x"833d0d04",
          6172 => x"fe3d0d76",
          6173 => x"75775454",
          6174 => x"5170802e",
          6175 => x"92387170",
          6176 => x"81055333",
          6177 => x"73708105",
          6178 => x"5534ff11",
          6179 => x"51eb3984",
          6180 => x"3d0d04fe",
          6181 => x"3d0d7577",
          6182 => x"76545253",
          6183 => x"72727081",
          6184 => x"055434ff",
          6185 => x"115170f4",
          6186 => x"38843d0d",
          6187 => x"04fc3d0d",
          6188 => x"78777956",
          6189 => x"56537470",
          6190 => x"81055633",
          6191 => x"74708105",
          6192 => x"56337171",
          6193 => x"31ff1656",
          6194 => x"52525272",
          6195 => x"802e8638",
          6196 => x"71802ee2",
          6197 => x"38718285",
          6198 => x"ec0c863d",
          6199 => x"0d04fe3d",
          6200 => x"0d747654",
          6201 => x"51893971",
          6202 => x"732e8a38",
          6203 => x"81115170",
          6204 => x"335271f3",
          6205 => x"38703382",
          6206 => x"85ec0c84",
          6207 => x"3d0d0480",
          6208 => x"0b8285ec",
          6209 => x"0c04800b",
          6210 => x"8285ec0c",
          6211 => x"04f73d0d",
          6212 => x"7b56800b",
          6213 => x"83173356",
          6214 => x"5a747a2e",
          6215 => x"80d63881",
          6216 => x"54b01608",
          6217 => x"53b41670",
          6218 => x"53811733",
          6219 => x"5259faa2",
          6220 => x"3f8285ec",
          6221 => x"087a2e09",
          6222 => x"8106b738",
          6223 => x"8285ec08",
          6224 => x"831734b0",
          6225 => x"160870a4",
          6226 => x"1808319c",
          6227 => x"18085956",
          6228 => x"58747727",
          6229 => x"9f388216",
          6230 => x"33557482",
          6231 => x"2e098106",
          6232 => x"93388154",
          6233 => x"76185378",
          6234 => x"52811633",
          6235 => x"51f9e33f",
          6236 => x"8339815a",
          6237 => x"798285ec",
          6238 => x"0c8b3d0d",
          6239 => x"04fa3d0d",
          6240 => x"787a5656",
          6241 => x"805774b0",
          6242 => x"17082eaf",
          6243 => x"387551fe",
          6244 => x"fc3f8285",
          6245 => x"ec085782",
          6246 => x"85ec089f",
          6247 => x"38815474",
          6248 => x"53b41652",
          6249 => x"81163351",
          6250 => x"f7be3f82",
          6251 => x"85ec0880",
          6252 => x"2e8538ff",
          6253 => x"55815774",
          6254 => x"b0170c76",
          6255 => x"8285ec0c",
          6256 => x"883d0d04",
          6257 => x"f83d0d7a",
          6258 => x"705257fe",
          6259 => x"c03f8285",
          6260 => x"ec085882",
          6261 => x"85ec0881",
          6262 => x"91387633",
          6263 => x"5574832e",
          6264 => x"09810680",
          6265 => x"f0388417",
          6266 => x"33597881",
          6267 => x"2e098106",
          6268 => x"80e33884",
          6269 => x"80538285",
          6270 => x"ec0852b4",
          6271 => x"17705256",
          6272 => x"fd913f82",
          6273 => x"d4d55284",
          6274 => x"b21751fc",
          6275 => x"963f848b",
          6276 => x"85a4d252",
          6277 => x"7551fca9",
          6278 => x"3f868a85",
          6279 => x"e4f25284",
          6280 => x"981751fc",
          6281 => x"9c3f9017",
          6282 => x"0852849c",
          6283 => x"1751fc91",
          6284 => x"3f8c1708",
          6285 => x"5284a017",
          6286 => x"51fc863f",
          6287 => x"a0170881",
          6288 => x"0570b019",
          6289 => x"0c795553",
          6290 => x"75528117",
          6291 => x"3351f882",
          6292 => x"3f778418",
          6293 => x"34805380",
          6294 => x"52811733",
          6295 => x"51f9d73f",
          6296 => x"8285ec08",
          6297 => x"802e8338",
          6298 => x"81587782",
          6299 => x"85ec0c8a",
          6300 => x"3d0d04fb",
          6301 => x"3d0d77fe",
          6302 => x"1a981208",
          6303 => x"fe055555",
          6304 => x"55805673",
          6305 => x"73279438",
          6306 => x"8a152274",
          6307 => x"5351ff97",
          6308 => x"f93fac15",
          6309 => x"088285ec",
          6310 => x"08055675",
          6311 => x"8285ec0c",
          6312 => x"873d0d04",
          6313 => x"f93d0d7a",
          6314 => x"7a700856",
          6315 => x"54578177",
          6316 => x"2781df38",
          6317 => x"76981508",
          6318 => x"2781d738",
          6319 => x"ff743354",
          6320 => x"5872822e",
          6321 => x"80f53872",
          6322 => x"82248938",
          6323 => x"72812e8d",
          6324 => x"3881bf39",
          6325 => x"72832e81",
          6326 => x"8e3881b6",
          6327 => x"3976812a",
          6328 => x"1770892a",
          6329 => x"a4160805",
          6330 => x"53745255",
          6331 => x"fd8f3f82",
          6332 => x"85ec0881",
          6333 => x"9f387483",
          6334 => x"ff0614b4",
          6335 => x"11338117",
          6336 => x"70892aa4",
          6337 => x"18080555",
          6338 => x"76545757",
          6339 => x"53fcee3f",
          6340 => x"8285ec08",
          6341 => x"80fe3874",
          6342 => x"83ff0614",
          6343 => x"b4113370",
          6344 => x"882b7807",
          6345 => x"79810671",
          6346 => x"842a5c52",
          6347 => x"58515372",
          6348 => x"80e23875",
          6349 => x"9fff0658",
          6350 => x"80da3976",
          6351 => x"882aa415",
          6352 => x"08055273",
          6353 => x"51fcb63f",
          6354 => x"8285ec08",
          6355 => x"80c63876",
          6356 => x"1083fe06",
          6357 => x"7405b405",
          6358 => x"51f9863f",
          6359 => x"8285ec08",
          6360 => x"83ffff06",
          6361 => x"58ae3976",
          6362 => x"872aa415",
          6363 => x"08055273",
          6364 => x"51fc8a3f",
          6365 => x"8285ec08",
          6366 => x"9b387682",
          6367 => x"2b83fc06",
          6368 => x"7405b405",
          6369 => x"51f8f13f",
          6370 => x"8285ec08",
          6371 => x"f00a0658",
          6372 => x"83398158",
          6373 => x"778285ec",
          6374 => x"0c893d0d",
          6375 => x"04f83d0d",
          6376 => x"7a7c7e5a",
          6377 => x"58568259",
          6378 => x"81772782",
          6379 => x"9e387698",
          6380 => x"17082782",
          6381 => x"96387533",
          6382 => x"5372792e",
          6383 => x"819d3872",
          6384 => x"79248938",
          6385 => x"72812e8d",
          6386 => x"38828039",
          6387 => x"72832e81",
          6388 => x"b83881f7",
          6389 => x"3976812a",
          6390 => x"1770892a",
          6391 => x"a4180805",
          6392 => x"53765255",
          6393 => x"fb973f82",
          6394 => x"85ec0859",
          6395 => x"8285ec08",
          6396 => x"81d93874",
          6397 => x"83ff0616",
          6398 => x"b4058116",
          6399 => x"78810659",
          6400 => x"56547753",
          6401 => x"76802e8f",
          6402 => x"3877842b",
          6403 => x"9ff00674",
          6404 => x"338f0671",
          6405 => x"07515372",
          6406 => x"7434810b",
          6407 => x"83173474",
          6408 => x"892aa417",
          6409 => x"08055275",
          6410 => x"51fad23f",
          6411 => x"8285ec08",
          6412 => x"598285ec",
          6413 => x"08819438",
          6414 => x"7483ff06",
          6415 => x"16b40578",
          6416 => x"842a5454",
          6417 => x"768f3877",
          6418 => x"882a7433",
          6419 => x"81f00671",
          6420 => x"8f060751",
          6421 => x"53727434",
          6422 => x"80ec3976",
          6423 => x"882aa417",
          6424 => x"08055275",
          6425 => x"51fa963f",
          6426 => x"8285ec08",
          6427 => x"598285ec",
          6428 => x"0880d838",
          6429 => x"7783ffff",
          6430 => x"06527610",
          6431 => x"83fe0676",
          6432 => x"05b40551",
          6433 => x"f79d3fbe",
          6434 => x"3976872a",
          6435 => x"a4170805",
          6436 => x"527551f9",
          6437 => x"e83f8285",
          6438 => x"ec085982",
          6439 => x"85ec08ab",
          6440 => x"3877f00a",
          6441 => x"0677822b",
          6442 => x"83fc0670",
          6443 => x"18b40570",
          6444 => x"54515454",
          6445 => x"f6c23f82",
          6446 => x"85ec088f",
          6447 => x"0a067407",
          6448 => x"527251f6",
          6449 => x"fc3f810b",
          6450 => x"83173478",
          6451 => x"8285ec0c",
          6452 => x"8a3d0d04",
          6453 => x"f83d0d7a",
          6454 => x"7c7e7208",
          6455 => x"59565659",
          6456 => x"817527a4",
          6457 => x"38749817",
          6458 => x"08279d38",
          6459 => x"73802eaa",
          6460 => x"38ff5373",
          6461 => x"527551fd",
          6462 => x"a43f8285",
          6463 => x"ec085482",
          6464 => x"85ec0880",
          6465 => x"f2389339",
          6466 => x"825480eb",
          6467 => x"39815480",
          6468 => x"e6398285",
          6469 => x"ec085480",
          6470 => x"de397452",
          6471 => x"7851fb84",
          6472 => x"3f8285ec",
          6473 => x"08588285",
          6474 => x"ec08802e",
          6475 => x"80c73882",
          6476 => x"85ec0881",
          6477 => x"2ed23882",
          6478 => x"85ec08ff",
          6479 => x"2ecf3880",
          6480 => x"53745275",
          6481 => x"51fcd63f",
          6482 => x"8285ec08",
          6483 => x"c5389816",
          6484 => x"08fe1190",
          6485 => x"18085755",
          6486 => x"57747427",
          6487 => x"90388115",
          6488 => x"90170c84",
          6489 => x"16338107",
          6490 => x"54738417",
          6491 => x"34775576",
          6492 => x"7826ffa6",
          6493 => x"38805473",
          6494 => x"8285ec0c",
          6495 => x"8a3d0d04",
          6496 => x"f63d0d7c",
          6497 => x"7e710859",
          6498 => x"5b5b7995",
          6499 => x"388c1708",
          6500 => x"5877802e",
          6501 => x"88389817",
          6502 => x"087826b2",
          6503 => x"388158ae",
          6504 => x"3979527a",
          6505 => x"51f9fd3f",
          6506 => x"81557482",
          6507 => x"85ec0827",
          6508 => x"82e63882",
          6509 => x"85ec0855",
          6510 => x"8285ec08",
          6511 => x"ff2e82d8",
          6512 => x"38981708",
          6513 => x"8285ec08",
          6514 => x"2682cd38",
          6515 => x"79589017",
          6516 => x"08705654",
          6517 => x"73802e82",
          6518 => x"bf38777a",
          6519 => x"2e098106",
          6520 => x"80e43881",
          6521 => x"1a569817",
          6522 => x"08762683",
          6523 => x"38825675",
          6524 => x"527a51f9",
          6525 => x"af3f8059",
          6526 => x"8285ec08",
          6527 => x"812e0981",
          6528 => x"06863882",
          6529 => x"85ec0859",
          6530 => x"8285ec08",
          6531 => x"09700981",
          6532 => x"05707207",
          6533 => x"8025707c",
          6534 => x"078285ec",
          6535 => x"08545151",
          6536 => x"55557381",
          6537 => x"f3388285",
          6538 => x"ec08802e",
          6539 => x"95388c17",
          6540 => x"08548174",
          6541 => x"27903873",
          6542 => x"98180827",
          6543 => x"89387358",
          6544 => x"85397580",
          6545 => x"dd387756",
          6546 => x"81165698",
          6547 => x"17087626",
          6548 => x"89388256",
          6549 => x"75782681",
          6550 => x"b0387552",
          6551 => x"7a51f8c4",
          6552 => x"3f8285ec",
          6553 => x"08802eba",
          6554 => x"38805982",
          6555 => x"85ec0881",
          6556 => x"2e098106",
          6557 => x"86388285",
          6558 => x"ec085982",
          6559 => x"85ec0809",
          6560 => x"70098105",
          6561 => x"70720780",
          6562 => x"25707c07",
          6563 => x"51515555",
          6564 => x"7380fa38",
          6565 => x"75782e09",
          6566 => x"8106ffac",
          6567 => x"38735580",
          6568 => x"f739ff53",
          6569 => x"75527651",
          6570 => x"f9f33f82",
          6571 => x"85ec0882",
          6572 => x"85ec0809",
          6573 => x"81057082",
          6574 => x"85ec0807",
          6575 => x"80255155",
          6576 => x"5579802e",
          6577 => x"94387380",
          6578 => x"2e8f3875",
          6579 => x"53795276",
          6580 => x"51f9ca3f",
          6581 => x"8285ec08",
          6582 => x"5574a538",
          6583 => x"758c180c",
          6584 => x"981708fe",
          6585 => x"05901808",
          6586 => x"56547474",
          6587 => x"268638ff",
          6588 => x"1590180c",
          6589 => x"84173381",
          6590 => x"07547384",
          6591 => x"18349739",
          6592 => x"ff567481",
          6593 => x"2e90388c",
          6594 => x"3980558c",
          6595 => x"398285ec",
          6596 => x"08558539",
          6597 => x"81567555",
          6598 => x"748285ec",
          6599 => x"0c8c3d0d",
          6600 => x"04f83d0d",
          6601 => x"7a705255",
          6602 => x"f3e33f82",
          6603 => x"85ec0858",
          6604 => x"81568285",
          6605 => x"ec0880da",
          6606 => x"387b5274",
          6607 => x"51f6b43f",
          6608 => x"8285ec08",
          6609 => x"8285ec08",
          6610 => x"b0170c59",
          6611 => x"84805377",
          6612 => x"52b41570",
          6613 => x"5257f2bb",
          6614 => x"3f775684",
          6615 => x"39811656",
          6616 => x"8a152258",
          6617 => x"75782797",
          6618 => x"38815475",
          6619 => x"19537652",
          6620 => x"81153351",
          6621 => x"eddc3f82",
          6622 => x"85ec0880",
          6623 => x"2edf388a",
          6624 => x"15227632",
          6625 => x"70098105",
          6626 => x"70720770",
          6627 => x"9f2a5351",
          6628 => x"56567582",
          6629 => x"85ec0c8a",
          6630 => x"3d0d04f8",
          6631 => x"3d0d7a7c",
          6632 => x"71085856",
          6633 => x"5774f080",
          6634 => x"0a2680f1",
          6635 => x"38749f06",
          6636 => x"537280e9",
          6637 => x"38749018",
          6638 => x"0c881708",
          6639 => x"5473aa38",
          6640 => x"75335382",
          6641 => x"73278838",
          6642 => x"a8160854",
          6643 => x"739b3874",
          6644 => x"852a5382",
          6645 => x"0b881722",
          6646 => x"5a587279",
          6647 => x"2780fe38",
          6648 => x"a8160898",
          6649 => x"180c80cd",
          6650 => x"398a1622",
          6651 => x"70892b54",
          6652 => x"58727526",
          6653 => x"b2387352",
          6654 => x"7651f5a8",
          6655 => x"3f8285ec",
          6656 => x"08548285",
          6657 => x"ec08ff2e",
          6658 => x"bd38810b",
          6659 => x"8285ec08",
          6660 => x"278b3898",
          6661 => x"16088285",
          6662 => x"ec082685",
          6663 => x"388258bd",
          6664 => x"39747331",
          6665 => x"55cb3973",
          6666 => x"527551f4",
          6667 => x"c63f8285",
          6668 => x"ec089818",
          6669 => x"0c739418",
          6670 => x"0c981708",
          6671 => x"53825872",
          6672 => x"802e9a38",
          6673 => x"85398158",
          6674 => x"94397489",
          6675 => x"2a139818",
          6676 => x"0c7483ff",
          6677 => x"0616b405",
          6678 => x"9c180c80",
          6679 => x"58778285",
          6680 => x"ec0c8a3d",
          6681 => x"0d04f83d",
          6682 => x"0d7a7008",
          6683 => x"901208a0",
          6684 => x"05595754",
          6685 => x"f0800a77",
          6686 => x"27863880",
          6687 => x"0b98150c",
          6688 => x"98140853",
          6689 => x"84557280",
          6690 => x"2e81cb38",
          6691 => x"7683ff06",
          6692 => x"587781b5",
          6693 => x"38811398",
          6694 => x"150c9414",
          6695 => x"08557492",
          6696 => x"3876852a",
          6697 => x"88172256",
          6698 => x"53747326",
          6699 => x"819b3880",
          6700 => x"c0398a16",
          6701 => x"22ff0577",
          6702 => x"892a0653",
          6703 => x"72818a38",
          6704 => x"74527351",
          6705 => x"f3de3f82",
          6706 => x"85ec0853",
          6707 => x"8255810b",
          6708 => x"8285ec08",
          6709 => x"2780ff38",
          6710 => x"81558285",
          6711 => x"ec08ff2e",
          6712 => x"80f43898",
          6713 => x"16088285",
          6714 => x"ec082680",
          6715 => x"ca387b8a",
          6716 => x"38779815",
          6717 => x"0c845580",
          6718 => x"dd399414",
          6719 => x"08527351",
          6720 => x"f8fe3f82",
          6721 => x"85ec0853",
          6722 => x"87558285",
          6723 => x"ec08802e",
          6724 => x"80c43882",
          6725 => x"558285ec",
          6726 => x"08812eba",
          6727 => x"38815582",
          6728 => x"85ec08ff",
          6729 => x"2eb03882",
          6730 => x"85ec0852",
          6731 => x"7551fbf1",
          6732 => x"3f8285ec",
          6733 => x"08a03872",
          6734 => x"94150c72",
          6735 => x"527551f2",
          6736 => x"b23f8285",
          6737 => x"ec089815",
          6738 => x"0c769015",
          6739 => x"0c7716b4",
          6740 => x"059c150c",
          6741 => x"80557482",
          6742 => x"85ec0c8a",
          6743 => x"3d0d04f7",
          6744 => x"3d0d7b7d",
          6745 => x"71085b5b",
          6746 => x"57805276",
          6747 => x"51fcac3f",
          6748 => x"8285ec08",
          6749 => x"548285ec",
          6750 => x"0880ec38",
          6751 => x"8285ec08",
          6752 => x"56981708",
          6753 => x"527851ef",
          6754 => x"f43f8285",
          6755 => x"ec085482",
          6756 => x"85ec0880",
          6757 => x"d2388285",
          6758 => x"ec089c18",
          6759 => x"08703351",
          6760 => x"54587281",
          6761 => x"e52e0981",
          6762 => x"06833881",
          6763 => x"588285ec",
          6764 => x"08557283",
          6765 => x"38815577",
          6766 => x"75075372",
          6767 => x"802e8e38",
          6768 => x"81165675",
          6769 => x"7a2e0981",
          6770 => x"068838a5",
          6771 => x"398285ec",
          6772 => x"08568152",
          6773 => x"7651fd8e",
          6774 => x"3f8285ec",
          6775 => x"08548285",
          6776 => x"ec08802e",
          6777 => x"ff9b3873",
          6778 => x"842e0981",
          6779 => x"06833887",
          6780 => x"54738285",
          6781 => x"ec0c8b3d",
          6782 => x"0d04fd3d",
          6783 => x"0d769a11",
          6784 => x"5254ebdd",
          6785 => x"3f8285ec",
          6786 => x"0883ffff",
          6787 => x"06767033",
          6788 => x"51535371",
          6789 => x"832e0981",
          6790 => x"06903894",
          6791 => x"1451ebc1",
          6792 => x"3f8285ec",
          6793 => x"08902b73",
          6794 => x"07537282",
          6795 => x"85ec0c85",
          6796 => x"3d0d04fc",
          6797 => x"3d0d7779",
          6798 => x"7083ffff",
          6799 => x"06549a12",
          6800 => x"535555eb",
          6801 => x"de3f7670",
          6802 => x"33515372",
          6803 => x"832e0981",
          6804 => x"068b3873",
          6805 => x"902a5294",
          6806 => x"1551ebc7",
          6807 => x"3f863d0d",
          6808 => x"04f73d0d",
          6809 => x"7b7d5b55",
          6810 => x"8475085a",
          6811 => x"58981508",
          6812 => x"802e818a",
          6813 => x"38981508",
          6814 => x"527851ee",
          6815 => x"803f8285",
          6816 => x"ec085882",
          6817 => x"85ec0880",
          6818 => x"f5389c15",
          6819 => x"08703355",
          6820 => x"53738638",
          6821 => x"845880e6",
          6822 => x"398b1333",
          6823 => x"70bf0670",
          6824 => x"81ff0658",
          6825 => x"51537286",
          6826 => x"16348285",
          6827 => x"ec085373",
          6828 => x"81e52e83",
          6829 => x"38815373",
          6830 => x"ae2ea938",
          6831 => x"81707406",
          6832 => x"54577280",
          6833 => x"2e9e3875",
          6834 => x"8f2e9938",
          6835 => x"8285ec08",
          6836 => x"76df0654",
          6837 => x"5472882e",
          6838 => x"09810683",
          6839 => x"38765473",
          6840 => x"7a2ea038",
          6841 => x"80527451",
          6842 => x"fafc3f82",
          6843 => x"85ec0858",
          6844 => x"8285ec08",
          6845 => x"89389815",
          6846 => x"08fefa38",
          6847 => x"8639800b",
          6848 => x"98160c77",
          6849 => x"8285ec0c",
          6850 => x"8b3d0d04",
          6851 => x"fb3d0d77",
          6852 => x"70085754",
          6853 => x"81527351",
          6854 => x"fcc53f82",
          6855 => x"85ec0855",
          6856 => x"8285ec08",
          6857 => x"b4389814",
          6858 => x"08527551",
          6859 => x"eccf3f82",
          6860 => x"85ec0855",
          6861 => x"8285ec08",
          6862 => x"a038a053",
          6863 => x"8285ec08",
          6864 => x"529c1408",
          6865 => x"51eacc3f",
          6866 => x"8b53a014",
          6867 => x"529c1408",
          6868 => x"51ea9d3f",
          6869 => x"810b8317",
          6870 => x"34748285",
          6871 => x"ec0c873d",
          6872 => x"0d04fd3d",
          6873 => x"0d757008",
          6874 => x"98120854",
          6875 => x"70535553",
          6876 => x"ec8b3f82",
          6877 => x"85ec088d",
          6878 => x"389c1308",
          6879 => x"53e57334",
          6880 => x"810b8315",
          6881 => x"34853d0d",
          6882 => x"04fa3d0d",
          6883 => x"787a5757",
          6884 => x"800b8917",
          6885 => x"34981708",
          6886 => x"802e8182",
          6887 => x"38807089",
          6888 => x"18555555",
          6889 => x"9c170814",
          6890 => x"70338116",
          6891 => x"56515271",
          6892 => x"a02ea838",
          6893 => x"71852e09",
          6894 => x"81068438",
          6895 => x"81e55273",
          6896 => x"892e0981",
          6897 => x"068b38ae",
          6898 => x"73708105",
          6899 => x"55348115",
          6900 => x"55717370",
          6901 => x"81055534",
          6902 => x"8115558a",
          6903 => x"7427c538",
          6904 => x"75158805",
          6905 => x"52800b81",
          6906 => x"13349c17",
          6907 => x"08528b12",
          6908 => x"33881734",
          6909 => x"9c17089c",
          6910 => x"115252e7",
          6911 => x"fb3f8285",
          6912 => x"ec08760c",
          6913 => x"961251e7",
          6914 => x"d83f8285",
          6915 => x"ec088617",
          6916 => x"23981251",
          6917 => x"e7cb3f82",
          6918 => x"85ec0884",
          6919 => x"1723883d",
          6920 => x"0d04f33d",
          6921 => x"0d7f7008",
          6922 => x"5e5b8061",
          6923 => x"70335155",
          6924 => x"5573af2e",
          6925 => x"83388155",
          6926 => x"7380dc2e",
          6927 => x"91387480",
          6928 => x"2e8c3894",
          6929 => x"1d08881c",
          6930 => x"0cac3981",
          6931 => x"15418061",
          6932 => x"70335656",
          6933 => x"5673af2e",
          6934 => x"09810683",
          6935 => x"38815673",
          6936 => x"80dc3270",
          6937 => x"09810570",
          6938 => x"80257807",
          6939 => x"51515473",
          6940 => x"da387388",
          6941 => x"1c0c6070",
          6942 => x"33515473",
          6943 => x"9f269638",
          6944 => x"ff800bab",
          6945 => x"1c348052",
          6946 => x"7a51f68f",
          6947 => x"3f8285ec",
          6948 => x"085585a6",
          6949 => x"39913d61",
          6950 => x"a01d5c5a",
          6951 => x"5e8b53a0",
          6952 => x"527951e7",
          6953 => x"ee3f8070",
          6954 => x"59578879",
          6955 => x"33555c73",
          6956 => x"ae2e0981",
          6957 => x"0680d838",
          6958 => x"78187033",
          6959 => x"811a71ae",
          6960 => x"32700981",
          6961 => x"05709f2a",
          6962 => x"73822607",
          6963 => x"5151535a",
          6964 => x"5754738c",
          6965 => x"38791754",
          6966 => x"75743481",
          6967 => x"1757d939",
          6968 => x"75af3270",
          6969 => x"09810570",
          6970 => x"9f2a5151",
          6971 => x"547580dc",
          6972 => x"2e8c3873",
          6973 => x"802e8738",
          6974 => x"75a02682",
          6975 => x"c7387719",
          6976 => x"7e0ca454",
          6977 => x"a0762782",
          6978 => x"c738a054",
          6979 => x"82c23978",
          6980 => x"18703381",
          6981 => x"1a5a5754",
          6982 => x"a0762782",
          6983 => x"863875af",
          6984 => x"32700981",
          6985 => x"057780dc",
          6986 => x"32700981",
          6987 => x"05728025",
          6988 => x"71802507",
          6989 => x"51515651",
          6990 => x"5573802e",
          6991 => x"ae388439",
          6992 => x"81185880",
          6993 => x"781a7033",
          6994 => x"51555573",
          6995 => x"af2e0981",
          6996 => x"06833881",
          6997 => x"557380dc",
          6998 => x"32700981",
          6999 => x"05708025",
          7000 => x"77075151",
          7001 => x"5473d938",
          7002 => x"81b93975",
          7003 => x"ae2e0981",
          7004 => x"06833881",
          7005 => x"54767c27",
          7006 => x"74075473",
          7007 => x"802ea638",
          7008 => x"7b8b3270",
          7009 => x"09810577",
          7010 => x"ae327009",
          7011 => x"81057280",
          7012 => x"25719f2a",
          7013 => x"07535156",
          7014 => x"51557481",
          7015 => x"a7388857",
          7016 => x"8b5cfeeb",
          7017 => x"3975982b",
          7018 => x"54738025",
          7019 => x"8c387580",
          7020 => x"ff0681ff",
          7021 => x"b4113357",
          7022 => x"547551e6",
          7023 => x"c23f8285",
          7024 => x"ec08802e",
          7025 => x"b2387818",
          7026 => x"7033811a",
          7027 => x"71545a56",
          7028 => x"54e6b33f",
          7029 => x"8285ec08",
          7030 => x"802e80e8",
          7031 => x"38ff1c54",
          7032 => x"76742780",
          7033 => x"df387917",
          7034 => x"54757434",
          7035 => x"81177a11",
          7036 => x"55577474",
          7037 => x"34a73975",
          7038 => x"5281fed4",
          7039 => x"51e5df3f",
          7040 => x"8285ec08",
          7041 => x"bf38ff9f",
          7042 => x"16547399",
          7043 => x"268938e0",
          7044 => x"167081ff",
          7045 => x"06575479",
          7046 => x"17547574",
          7047 => x"34811757",
          7048 => x"fded3977",
          7049 => x"197e0c76",
          7050 => x"802e9938",
          7051 => x"79335473",
          7052 => x"81e52e09",
          7053 => x"81068438",
          7054 => x"857a3484",
          7055 => x"54a07627",
          7056 => x"8f388b39",
          7057 => x"865581f2",
          7058 => x"39845680",
          7059 => x"f3398054",
          7060 => x"738b1b34",
          7061 => x"807b0858",
          7062 => x"527a51f2",
          7063 => x"be3f8285",
          7064 => x"ec085682",
          7065 => x"85ec0880",
          7066 => x"d738981b",
          7067 => x"08527651",
          7068 => x"e68b3f82",
          7069 => x"85ec0856",
          7070 => x"8285ec08",
          7071 => x"80c2389c",
          7072 => x"1b087033",
          7073 => x"55557380",
          7074 => x"2effbe38",
          7075 => x"8b1533bf",
          7076 => x"06547386",
          7077 => x"1c348b15",
          7078 => x"3370832a",
          7079 => x"70810651",
          7080 => x"55587392",
          7081 => x"388b5379",
          7082 => x"527451e4",
          7083 => x"803f8285",
          7084 => x"ec08802e",
          7085 => x"8b387552",
          7086 => x"7a51f3aa",
          7087 => x"3fff9f39",
          7088 => x"75ab1c33",
          7089 => x"57557480",
          7090 => x"2ebb3874",
          7091 => x"842e0981",
          7092 => x"0680e738",
          7093 => x"75852a70",
          7094 => x"81067782",
          7095 => x"2a585154",
          7096 => x"73802e96",
          7097 => x"38758106",
          7098 => x"5473802e",
          7099 => x"fba738ff",
          7100 => x"800bab1c",
          7101 => x"34805580",
          7102 => x"c1397581",
          7103 => x"065473ba",
          7104 => x"388555b6",
          7105 => x"3975822a",
          7106 => x"70810651",
          7107 => x"5473ab38",
          7108 => x"861b3370",
          7109 => x"842a7081",
          7110 => x"06515555",
          7111 => x"73802ee1",
          7112 => x"38901b08",
          7113 => x"83ff061d",
          7114 => x"b405527c",
          7115 => x"51f5cb3f",
          7116 => x"8285ec08",
          7117 => x"881c0cfa",
          7118 => x"dc397482",
          7119 => x"85ec0c8f",
          7120 => x"3d0d04f6",
          7121 => x"3d0d7c5b",
          7122 => x"ff7b0870",
          7123 => x"71735559",
          7124 => x"5c555973",
          7125 => x"802e81cc",
          7126 => x"38757081",
          7127 => x"05573370",
          7128 => x"a0265252",
          7129 => x"71ba2e8d",
          7130 => x"3870ee38",
          7131 => x"71ba2e09",
          7132 => x"810681ab",
          7133 => x"387333d0",
          7134 => x"117081ff",
          7135 => x"06515253",
          7136 => x"70892691",
          7137 => x"38821473",
          7138 => x"81ff06d0",
          7139 => x"05565271",
          7140 => x"762e80fd",
          7141 => x"38800b81",
          7142 => x"ffa45955",
          7143 => x"77087a55",
          7144 => x"57767081",
          7145 => x"05583374",
          7146 => x"70810556",
          7147 => x"33ff9f12",
          7148 => x"53535370",
          7149 => x"99268938",
          7150 => x"e0137081",
          7151 => x"ff065451",
          7152 => x"ff9f1251",
          7153 => x"70992689",
          7154 => x"38e01270",
          7155 => x"81ff0653",
          7156 => x"51720981",
          7157 => x"05709f2a",
          7158 => x"51517272",
          7159 => x"2e098106",
          7160 => x"853870ff",
          7161 => x"bc387209",
          7162 => x"81057477",
          7163 => x"32700981",
          7164 => x"05707207",
          7165 => x"9f2a739f",
          7166 => x"2a075354",
          7167 => x"54517080",
          7168 => x"2e8f3881",
          7169 => x"15841959",
          7170 => x"55837525",
          7171 => x"ff8e388b",
          7172 => x"39748324",
          7173 => x"86387476",
          7174 => x"7c0c5978",
          7175 => x"51863982",
          7176 => x"9da43351",
          7177 => x"708285ec",
          7178 => x"0c8c3d0d",
          7179 => x"04fa3d0d",
          7180 => x"7856800b",
          7181 => x"831734ff",
          7182 => x"0bb0170c",
          7183 => x"79527551",
          7184 => x"e2bb3f84",
          7185 => x"558285ec",
          7186 => x"08818238",
          7187 => x"84b21651",
          7188 => x"df8f3f82",
          7189 => x"85ec0883",
          7190 => x"ffff0654",
          7191 => x"83557382",
          7192 => x"d4d52e09",
          7193 => x"810680e5",
          7194 => x"38800bb4",
          7195 => x"17335657",
          7196 => x"7481e92e",
          7197 => x"09810683",
          7198 => x"38815774",
          7199 => x"81eb3270",
          7200 => x"09810570",
          7201 => x"80257907",
          7202 => x"51515473",
          7203 => x"8a387481",
          7204 => x"e82e0981",
          7205 => x"06b53883",
          7206 => x"5381fee4",
          7207 => x"5280ea16",
          7208 => x"51e08a3f",
          7209 => x"8285ec08",
          7210 => x"558285ec",
          7211 => x"08802e9d",
          7212 => x"38855381",
          7213 => x"fee85281",
          7214 => x"861651df",
          7215 => x"f03f8285",
          7216 => x"ec085582",
          7217 => x"85ec0880",
          7218 => x"2e833882",
          7219 => x"55748285",
          7220 => x"ec0c883d",
          7221 => x"0d04f13d",
          7222 => x"0d620284",
          7223 => x"0580cf05",
          7224 => x"33585580",
          7225 => x"750c6151",
          7226 => x"fcd93f82",
          7227 => x"85ec0858",
          7228 => x"8b56800b",
          7229 => x"8285ec08",
          7230 => x"24878338",
          7231 => x"8285ec08",
          7232 => x"822b829d",
          7233 => x"90110855",
          7234 => x"538c5673",
          7235 => x"802e86ee",
          7236 => x"3873750c",
          7237 => x"7681fe06",
          7238 => x"74335457",
          7239 => x"72802eae",
          7240 => x"38811433",
          7241 => x"51d7a43f",
          7242 => x"8285ec08",
          7243 => x"81ff0670",
          7244 => x"81065455",
          7245 => x"72983876",
          7246 => x"802e86c0",
          7247 => x"3874822a",
          7248 => x"70810651",
          7249 => x"538a5672",
          7250 => x"86b43886",
          7251 => x"af398074",
          7252 => x"34778115",
          7253 => x"34815281",
          7254 => x"143351d7",
          7255 => x"8c3f8285",
          7256 => x"ec0881ff",
          7257 => x"06708106",
          7258 => x"54558356",
          7259 => x"72868f38",
          7260 => x"76802e8f",
          7261 => x"3874822a",
          7262 => x"70810651",
          7263 => x"538a5672",
          7264 => x"85fc3880",
          7265 => x"70537452",
          7266 => x"5cfda23f",
          7267 => x"8285ec08",
          7268 => x"81ff0657",
          7269 => x"76822e09",
          7270 => x"810680e2",
          7271 => x"388d3d74",
          7272 => x"56588356",
          7273 => x"83f61533",
          7274 => x"70585372",
          7275 => x"802e8d38",
          7276 => x"83fa1551",
          7277 => x"dcc23f82",
          7278 => x"85ec0857",
          7279 => x"76787084",
          7280 => x"055a0cff",
          7281 => x"16901656",
          7282 => x"56758025",
          7283 => x"d738800b",
          7284 => x"8e3d5456",
          7285 => x"72708405",
          7286 => x"54085c83",
          7287 => x"577b802e",
          7288 => x"95387b52",
          7289 => x"7351fcc5",
          7290 => x"3f8285ec",
          7291 => x"0881ff06",
          7292 => x"57817727",
          7293 => x"89388116",
          7294 => x"56837627",
          7295 => x"d7388156",
          7296 => x"76842e84",
          7297 => x"f9388d56",
          7298 => x"76812684",
          7299 => x"f138bf14",
          7300 => x"51dbce3f",
          7301 => x"8285ec08",
          7302 => x"83ffff06",
          7303 => x"53728480",
          7304 => x"2e098106",
          7305 => x"84d83880",
          7306 => x"ca1451db",
          7307 => x"b43f8285",
          7308 => x"ec0883ff",
          7309 => x"ff065877",
          7310 => x"8d3880d8",
          7311 => x"1451dbb8",
          7312 => x"3f8285ec",
          7313 => x"0858779c",
          7314 => x"150c80c4",
          7315 => x"14338215",
          7316 => x"3480c414",
          7317 => x"33ff1170",
          7318 => x"81ff0651",
          7319 => x"54558d56",
          7320 => x"72812684",
          7321 => x"99387481",
          7322 => x"ff065277",
          7323 => x"51fef89a",
          7324 => x"3f8285ec",
          7325 => x"0880c115",
          7326 => x"33545872",
          7327 => x"8a152372",
          7328 => x"802e8b38",
          7329 => x"ff137306",
          7330 => x"5372802e",
          7331 => x"86388d56",
          7332 => x"83ec3980",
          7333 => x"c51451da",
          7334 => x"c83f8285",
          7335 => x"ec085382",
          7336 => x"85ec0888",
          7337 => x"1523728f",
          7338 => x"06578d56",
          7339 => x"7683cf38",
          7340 => x"80c71451",
          7341 => x"daab3f82",
          7342 => x"85ec0883",
          7343 => x"ffff0655",
          7344 => x"748d3880",
          7345 => x"d41451da",
          7346 => x"af3f8285",
          7347 => x"ec085580",
          7348 => x"c21451da",
          7349 => x"8c3f8285",
          7350 => x"ec0883ff",
          7351 => x"ff065a8d",
          7352 => x"5679802e",
          7353 => x"83983888",
          7354 => x"1422781b",
          7355 => x"71842a05",
          7356 => x"5a5b7875",
          7357 => x"26838738",
          7358 => x"8a142252",
          7359 => x"74793151",
          7360 => x"fef8873f",
          7361 => x"8285ec08",
          7362 => x"538285ec",
          7363 => x"08802e82",
          7364 => x"ed388285",
          7365 => x"ec0880ff",
          7366 => x"fffff526",
          7367 => x"83388357",
          7368 => x"7283fff5",
          7369 => x"26833882",
          7370 => x"57729ff5",
          7371 => x"26853881",
          7372 => x"5789398d",
          7373 => x"5676802e",
          7374 => x"82c43882",
          7375 => x"13709816",
          7376 => x"0c7ca016",
          7377 => x"0c7a1d70",
          7378 => x"a4170c7a",
          7379 => x"1eac170c",
          7380 => x"54557683",
          7381 => x"2e098106",
          7382 => x"af3880de",
          7383 => x"1451d981",
          7384 => x"3f8285ec",
          7385 => x"0883ffff",
          7386 => x"06538d56",
          7387 => x"72828f38",
          7388 => x"7a828b38",
          7389 => x"80e01451",
          7390 => x"d8fe3f82",
          7391 => x"85ec08a8",
          7392 => x"150c7482",
          7393 => x"2b53a339",
          7394 => x"8d567a80",
          7395 => x"2e81ef38",
          7396 => x"7713a815",
          7397 => x"0c741553",
          7398 => x"76822e8e",
          7399 => x"38741075",
          7400 => x"11812a76",
          7401 => x"81061151",
          7402 => x"515383ff",
          7403 => x"13892a53",
          7404 => x"8d56729c",
          7405 => x"15082681",
          7406 => x"c538ff0b",
          7407 => x"90150cff",
          7408 => x"0b8c150c",
          7409 => x"ff800b84",
          7410 => x"15347683",
          7411 => x"2e098106",
          7412 => x"81923880",
          7413 => x"e41451d8",
          7414 => x"883f8285",
          7415 => x"ec0883ff",
          7416 => x"ff065372",
          7417 => x"812e0981",
          7418 => x"0680f938",
          7419 => x"811c5273",
          7420 => x"51db8a3f",
          7421 => x"8285ec08",
          7422 => x"80ea3882",
          7423 => x"85ec0884",
          7424 => x"153484b2",
          7425 => x"1451d7d9",
          7426 => x"3f8285ec",
          7427 => x"0883ffff",
          7428 => x"06537282",
          7429 => x"d4d52e09",
          7430 => x"810680c8",
          7431 => x"38b41451",
          7432 => x"d7d63f82",
          7433 => x"85ec0884",
          7434 => x"8b85a4d2",
          7435 => x"2e098106",
          7436 => x"b3388498",
          7437 => x"1451d7c0",
          7438 => x"3f8285ec",
          7439 => x"08868a85",
          7440 => x"e4f22e09",
          7441 => x"81069d38",
          7442 => x"849c1451",
          7443 => x"d7aa3f82",
          7444 => x"85ec0890",
          7445 => x"150c84a0",
          7446 => x"1451d79c",
          7447 => x"3f8285ec",
          7448 => x"088c150c",
          7449 => x"76743482",
          7450 => x"9da02281",
          7451 => x"05537282",
          7452 => x"9da02372",
          7453 => x"86152380",
          7454 => x"0b94150c",
          7455 => x"80567582",
          7456 => x"85ec0c91",
          7457 => x"3d0d04fb",
          7458 => x"3d0d7754",
          7459 => x"89557380",
          7460 => x"2eb93873",
          7461 => x"08537280",
          7462 => x"2eb13872",
          7463 => x"33527180",
          7464 => x"2ea93886",
          7465 => x"13228415",
          7466 => x"22575271",
          7467 => x"762e0981",
          7468 => x"06993881",
          7469 => x"133351d0",
          7470 => x"923f8285",
          7471 => x"ec088106",
          7472 => x"52718838",
          7473 => x"71740854",
          7474 => x"55833980",
          7475 => x"53787371",
          7476 => x"0c527482",
          7477 => x"85ec0c87",
          7478 => x"3d0d04fa",
          7479 => x"3d0d02ab",
          7480 => x"05337a58",
          7481 => x"893dfc05",
          7482 => x"5256f4d7",
          7483 => x"3f8b5480",
          7484 => x"0b8285ec",
          7485 => x"0824bc38",
          7486 => x"8285ec08",
          7487 => x"822b829d",
          7488 => x"90057008",
          7489 => x"55557380",
          7490 => x"2e843880",
          7491 => x"74347854",
          7492 => x"73802e84",
          7493 => x"38807434",
          7494 => x"78750c75",
          7495 => x"5475802e",
          7496 => x"92388053",
          7497 => x"893d7053",
          7498 => x"840551f7",
          7499 => x"a93f8285",
          7500 => x"ec085473",
          7501 => x"8285ec0c",
          7502 => x"883d0d04",
          7503 => x"eb3d0d67",
          7504 => x"02840580",
          7505 => x"e7053359",
          7506 => x"59895478",
          7507 => x"802e84ca",
          7508 => x"3877bf06",
          7509 => x"7054983d",
          7510 => x"d0055399",
          7511 => x"3d840552",
          7512 => x"58f6f33f",
          7513 => x"8285ec08",
          7514 => x"558285ec",
          7515 => x"0884a638",
          7516 => x"7a5c6852",
          7517 => x"8c3d7052",
          7518 => x"56eda73f",
          7519 => x"8285ec08",
          7520 => x"558285ec",
          7521 => x"08923802",
          7522 => x"80d70533",
          7523 => x"70982b55",
          7524 => x"57738025",
          7525 => x"83388655",
          7526 => x"779c0654",
          7527 => x"73802e81",
          7528 => x"ab387480",
          7529 => x"2e953874",
          7530 => x"842e0981",
          7531 => x"06aa3875",
          7532 => x"51ead93f",
          7533 => x"8285ec08",
          7534 => x"559e3902",
          7535 => x"b2053391",
          7536 => x"06547381",
          7537 => x"b8387782",
          7538 => x"2a708106",
          7539 => x"51547380",
          7540 => x"2e8e3888",
          7541 => x"5583be39",
          7542 => x"77880758",
          7543 => x"7483b638",
          7544 => x"77832a70",
          7545 => x"81065154",
          7546 => x"73802e81",
          7547 => x"af386252",
          7548 => x"7a51e886",
          7549 => x"3f8285ec",
          7550 => x"08568288",
          7551 => x"b20a5262",
          7552 => x"8e0551d4",
          7553 => x"bc3f6254",
          7554 => x"a00b8b15",
          7555 => x"34805362",
          7556 => x"527a51e8",
          7557 => x"9e3f8052",
          7558 => x"629c0551",
          7559 => x"d4a33f7a",
          7560 => x"54810b83",
          7561 => x"15347580",
          7562 => x"2e80f138",
          7563 => x"7ab01108",
          7564 => x"51548053",
          7565 => x"7552973d",
          7566 => x"d40551dd",
          7567 => x"973f8285",
          7568 => x"ec085582",
          7569 => x"85ec0882",
          7570 => x"cc38b739",
          7571 => x"7482c638",
          7572 => x"02b20533",
          7573 => x"70842a70",
          7574 => x"81065155",
          7575 => x"5673802e",
          7576 => x"86388455",
          7577 => x"82af3977",
          7578 => x"812a7081",
          7579 => x"06515473",
          7580 => x"802ea938",
          7581 => x"75810654",
          7582 => x"73802ea0",
          7583 => x"38875582",
          7584 => x"94397352",
          7585 => x"7a51d5f5",
          7586 => x"3f8285ec",
          7587 => x"087bff18",
          7588 => x"8c120c55",
          7589 => x"558285ec",
          7590 => x"0881fa38",
          7591 => x"77832a70",
          7592 => x"81065154",
          7593 => x"73802e86",
          7594 => x"387780c0",
          7595 => x"07587ab0",
          7596 => x"1108a01b",
          7597 => x"0c63a41b",
          7598 => x"0c635370",
          7599 => x"5257e6ba",
          7600 => x"3f8285ec",
          7601 => x"088285ec",
          7602 => x"08881b0c",
          7603 => x"639c0552",
          7604 => x"5ad2a53f",
          7605 => x"8285ec08",
          7606 => x"8285ec08",
          7607 => x"8c1b0c77",
          7608 => x"7a0c5686",
          7609 => x"1722841a",
          7610 => x"2377901a",
          7611 => x"34800b91",
          7612 => x"1a34800b",
          7613 => x"9c1a0c80",
          7614 => x"0b941a0c",
          7615 => x"77852a70",
          7616 => x"81065154",
          7617 => x"73802e81",
          7618 => x"8f388285",
          7619 => x"ec08802e",
          7620 => x"81863882",
          7621 => x"85ec0894",
          7622 => x"1a0c8a17",
          7623 => x"2270892b",
          7624 => x"7b525957",
          7625 => x"a8397652",
          7626 => x"7851d6f8",
          7627 => x"3f8285ec",
          7628 => x"08578285",
          7629 => x"ec088126",
          7630 => x"83388255",
          7631 => x"8285ec08",
          7632 => x"ff2e0981",
          7633 => x"06833879",
          7634 => x"55757831",
          7635 => x"56740981",
          7636 => x"05707607",
          7637 => x"80255154",
          7638 => x"7776278a",
          7639 => x"38817075",
          7640 => x"06555a73",
          7641 => x"c1387698",
          7642 => x"1a0c74a9",
          7643 => x"387583ff",
          7644 => x"06547380",
          7645 => x"2ea23876",
          7646 => x"527a51d5",
          7647 => x"f63f8285",
          7648 => x"ec088538",
          7649 => x"82558e39",
          7650 => x"75892a82",
          7651 => x"85ec0805",
          7652 => x"9c1a0c84",
          7653 => x"3980790c",
          7654 => x"74547382",
          7655 => x"85ec0c97",
          7656 => x"3d0d04f2",
          7657 => x"3d0d6063",
          7658 => x"65644040",
          7659 => x"5d59807e",
          7660 => x"0c903dfc",
          7661 => x"05527851",
          7662 => x"f9cd3f82",
          7663 => x"85ec0855",
          7664 => x"8285ec08",
          7665 => x"8a389119",
          7666 => x"33557480",
          7667 => x"2e863874",
          7668 => x"5682c439",
          7669 => x"90193381",
          7670 => x"06558756",
          7671 => x"74802e82",
          7672 => x"b6389539",
          7673 => x"820b911a",
          7674 => x"34825682",
          7675 => x"aa39810b",
          7676 => x"911a3481",
          7677 => x"5682a039",
          7678 => x"8c190894",
          7679 => x"1a083155",
          7680 => x"747c2783",
          7681 => x"38745c7b",
          7682 => x"802e8289",
          7683 => x"38941908",
          7684 => x"7083ff06",
          7685 => x"56567481",
          7686 => x"b2387e8a",
          7687 => x"1122ff05",
          7688 => x"77892a06",
          7689 => x"5b5579a8",
          7690 => x"38758738",
          7691 => x"88190855",
          7692 => x"8f399819",
          7693 => x"08527851",
          7694 => x"d4ea3f82",
          7695 => x"85ec0855",
          7696 => x"817527ff",
          7697 => x"9f3874ff",
          7698 => x"2effa338",
          7699 => x"74981a0c",
          7700 => x"98190852",
          7701 => x"7e51d49b",
          7702 => x"3f8285ec",
          7703 => x"08802eff",
          7704 => x"83388285",
          7705 => x"ec081a7c",
          7706 => x"892a5957",
          7707 => x"77802e80",
          7708 => x"d638771a",
          7709 => x"7f8a1122",
          7710 => x"585c5575",
          7711 => x"75278538",
          7712 => x"757a3158",
          7713 => x"77547653",
          7714 => x"7c52811b",
          7715 => x"3351c9d8",
          7716 => x"3f8285ec",
          7717 => x"08fed738",
          7718 => x"7e831133",
          7719 => x"56567480",
          7720 => x"2e9f38b0",
          7721 => x"16087731",
          7722 => x"55747827",
          7723 => x"94388480",
          7724 => x"53b41652",
          7725 => x"b0160877",
          7726 => x"31892b7d",
          7727 => x"0551cfb0",
          7728 => x"3f77892b",
          7729 => x"56b93976",
          7730 => x"9c1a0c94",
          7731 => x"190883ff",
          7732 => x"06848071",
          7733 => x"3157557b",
          7734 => x"76278338",
          7735 => x"7b569c19",
          7736 => x"08527e51",
          7737 => x"d1973f82",
          7738 => x"85ec08fe",
          7739 => x"81387553",
          7740 => x"94190883",
          7741 => x"ff061fb4",
          7742 => x"05527c51",
          7743 => x"cef23f7b",
          7744 => x"76317e08",
          7745 => x"177f0c76",
          7746 => x"1e941b08",
          7747 => x"18941c0c",
          7748 => x"5e5cfdf3",
          7749 => x"39805675",
          7750 => x"8285ec0c",
          7751 => x"903d0d04",
          7752 => x"f23d0d60",
          7753 => x"63656440",
          7754 => x"405d5880",
          7755 => x"7e0c903d",
          7756 => x"fc055277",
          7757 => x"51f6d03f",
          7758 => x"8285ec08",
          7759 => x"558285ec",
          7760 => x"088a3891",
          7761 => x"18335574",
          7762 => x"802e8638",
          7763 => x"745683b8",
          7764 => x"39901833",
          7765 => x"70812a70",
          7766 => x"81065156",
          7767 => x"56875674",
          7768 => x"802e83a4",
          7769 => x"38953982",
          7770 => x"0b911934",
          7771 => x"82568398",
          7772 => x"39810b91",
          7773 => x"19348156",
          7774 => x"838e3994",
          7775 => x"18087c11",
          7776 => x"56567476",
          7777 => x"27843875",
          7778 => x"095c7b80",
          7779 => x"2e82ec38",
          7780 => x"94180870",
          7781 => x"83ff0656",
          7782 => x"567481fd",
          7783 => x"387e8a11",
          7784 => x"22ff0577",
          7785 => x"892a065c",
          7786 => x"557abf38",
          7787 => x"758c3888",
          7788 => x"18085574",
          7789 => x"9c387a52",
          7790 => x"85399818",
          7791 => x"08527751",
          7792 => x"d7be3f82",
          7793 => x"85ec0855",
          7794 => x"8285ec08",
          7795 => x"802e82ab",
          7796 => x"3874812e",
          7797 => x"ff913874",
          7798 => x"ff2eff95",
          7799 => x"38749819",
          7800 => x"0c881808",
          7801 => x"85387488",
          7802 => x"190c7e55",
          7803 => x"b015089c",
          7804 => x"19082e09",
          7805 => x"81068d38",
          7806 => x"7451ce91",
          7807 => x"3f8285ec",
          7808 => x"08feee38",
          7809 => x"98180852",
          7810 => x"7e51d0e7",
          7811 => x"3f8285ec",
          7812 => x"08802efe",
          7813 => x"d2388285",
          7814 => x"ec081b7c",
          7815 => x"892a5a57",
          7816 => x"78802e80",
          7817 => x"d538781b",
          7818 => x"7f8a1122",
          7819 => x"585b5575",
          7820 => x"75278538",
          7821 => x"757b3159",
          7822 => x"78547653",
          7823 => x"7c52811a",
          7824 => x"3351c88e",
          7825 => x"3f8285ec",
          7826 => x"08fea638",
          7827 => x"7eb01108",
          7828 => x"78315656",
          7829 => x"7479279b",
          7830 => x"38848053",
          7831 => x"b0160877",
          7832 => x"31892b7d",
          7833 => x"0552b416",
          7834 => x"51cc853f",
          7835 => x"7e55800b",
          7836 => x"83163478",
          7837 => x"892b5680",
          7838 => x"db398c18",
          7839 => x"08941908",
          7840 => x"2693387e",
          7841 => x"51cd863f",
          7842 => x"8285ec08",
          7843 => x"fde3387e",
          7844 => x"77b0120c",
          7845 => x"55769c19",
          7846 => x"0c941808",
          7847 => x"83ff0684",
          7848 => x"80713157",
          7849 => x"557b7627",
          7850 => x"83387b56",
          7851 => x"9c180852",
          7852 => x"7e51cdc9",
          7853 => x"3f8285ec",
          7854 => x"08fdb638",
          7855 => x"75537c52",
          7856 => x"94180883",
          7857 => x"ff061fb4",
          7858 => x"0551cba4",
          7859 => x"3f7e5581",
          7860 => x"0b831634",
          7861 => x"7b76317e",
          7862 => x"08177f0c",
          7863 => x"761e941a",
          7864 => x"08187094",
          7865 => x"1c0c8c1b",
          7866 => x"0858585e",
          7867 => x"5c747627",
          7868 => x"83387555",
          7869 => x"748c190c",
          7870 => x"fd903990",
          7871 => x"183380c0",
          7872 => x"07557490",
          7873 => x"19348056",
          7874 => x"758285ec",
          7875 => x"0c903d0d",
          7876 => x"04f83d0d",
          7877 => x"7a8b3dfc",
          7878 => x"05537052",
          7879 => x"56f2e83f",
          7880 => x"8285ec08",
          7881 => x"578285ec",
          7882 => x"0880fb38",
          7883 => x"90163370",
          7884 => x"862a7081",
          7885 => x"06515555",
          7886 => x"73802e80",
          7887 => x"e938a016",
          7888 => x"08527851",
          7889 => x"ccb73f82",
          7890 => x"85ec0857",
          7891 => x"8285ec08",
          7892 => x"80d438a4",
          7893 => x"16088b11",
          7894 => x"33a00755",
          7895 => x"55738b16",
          7896 => x"34881608",
          7897 => x"53745275",
          7898 => x"0851ddc7",
          7899 => x"3f8c1608",
          7900 => x"529c1551",
          7901 => x"c9cb3f82",
          7902 => x"88b20a52",
          7903 => x"961551c9",
          7904 => x"c03f7652",
          7905 => x"921551c9",
          7906 => x"9a3f7854",
          7907 => x"810b8315",
          7908 => x"347851cc",
          7909 => x"af3f8285",
          7910 => x"ec089017",
          7911 => x"3381bf06",
          7912 => x"55577390",
          7913 => x"17347682",
          7914 => x"85ec0c8a",
          7915 => x"3d0d04fc",
          7916 => x"3d0d7670",
          7917 => x"5254fed9",
          7918 => x"3f8285ec",
          7919 => x"08538285",
          7920 => x"ec089c38",
          7921 => x"863dfc05",
          7922 => x"527351f1",
          7923 => x"ba3f8285",
          7924 => x"ec085382",
          7925 => x"85ec0887",
          7926 => x"388285ec",
          7927 => x"08740c72",
          7928 => x"8285ec0c",
          7929 => x"863d0d04",
          7930 => x"ff3d0d84",
          7931 => x"3d51e6d3",
          7932 => x"3f8b5280",
          7933 => x"0b8285ec",
          7934 => x"08248b38",
          7935 => x"8285ec08",
          7936 => x"829da434",
          7937 => x"80527182",
          7938 => x"85ec0c83",
          7939 => x"3d0d04ef",
          7940 => x"3d0d8053",
          7941 => x"933dd005",
          7942 => x"52943d51",
          7943 => x"e9b83f82",
          7944 => x"85ec0855",
          7945 => x"8285ec08",
          7946 => x"80e03876",
          7947 => x"58635293",
          7948 => x"3dd40551",
          7949 => x"dfec3f82",
          7950 => x"85ec0855",
          7951 => x"8285ec08",
          7952 => x"bc380280",
          7953 => x"c7053370",
          7954 => x"982b5556",
          7955 => x"73802589",
          7956 => x"38767a94",
          7957 => x"120c54b2",
          7958 => x"3902a205",
          7959 => x"3370842a",
          7960 => x"70810651",
          7961 => x"55567380",
          7962 => x"2e9e3876",
          7963 => x"7f537052",
          7964 => x"54db873f",
          7965 => x"8285ec08",
          7966 => x"94150c8e",
          7967 => x"398285ec",
          7968 => x"08842e09",
          7969 => x"81068338",
          7970 => x"85557482",
          7971 => x"85ec0c93",
          7972 => x"3d0d04e4",
          7973 => x"3d0d6f6f",
          7974 => x"5b5b807a",
          7975 => x"3480539e",
          7976 => x"3dffb805",
          7977 => x"529f3d51",
          7978 => x"e8ac3f82",
          7979 => x"85ec0857",
          7980 => x"8285ec08",
          7981 => x"82fb387b",
          7982 => x"437a7c94",
          7983 => x"11084755",
          7984 => x"58645473",
          7985 => x"802e81ed",
          7986 => x"38a05293",
          7987 => x"3d705255",
          7988 => x"d5c93f82",
          7989 => x"85ec0857",
          7990 => x"8285ec08",
          7991 => x"82d33868",
          7992 => x"527b51c9",
          7993 => x"983f8285",
          7994 => x"ec085782",
          7995 => x"85ec0882",
          7996 => x"c0386952",
          7997 => x"7b51da82",
          7998 => x"3f8285ec",
          7999 => x"08457652",
          8000 => x"7451d597",
          8001 => x"3f8285ec",
          8002 => x"08578285",
          8003 => x"ec0882a1",
          8004 => x"38805274",
          8005 => x"51daca3f",
          8006 => x"8285ec08",
          8007 => x"578285ec",
          8008 => x"08a43869",
          8009 => x"527b51d9",
          8010 => x"d13f7382",
          8011 => x"85ec082e",
          8012 => x"a6387652",
          8013 => x"7451d6ae",
          8014 => x"3f8285ec",
          8015 => x"08578285",
          8016 => x"ec08802e",
          8017 => x"cc387684",
          8018 => x"2e098106",
          8019 => x"86388257",
          8020 => x"81df3976",
          8021 => x"81db389e",
          8022 => x"3dffbc05",
          8023 => x"527451dc",
          8024 => x"a83f7690",
          8025 => x"3d781181",
          8026 => x"11335156",
          8027 => x"5a567380",
          8028 => x"2e913802",
          8029 => x"b9055581",
          8030 => x"16811670",
          8031 => x"33565656",
          8032 => x"73f53881",
          8033 => x"16547378",
          8034 => x"26818f38",
          8035 => x"75802e99",
          8036 => x"38781681",
          8037 => x"0555ff18",
          8038 => x"6f11ff18",
          8039 => x"ff185858",
          8040 => x"55587433",
          8041 => x"743475ee",
          8042 => x"38ff186f",
          8043 => x"115558af",
          8044 => x"7434fe8d",
          8045 => x"39777b2e",
          8046 => x"0981068a",
          8047 => x"38ff186f",
          8048 => x"115558af",
          8049 => x"7434800b",
          8050 => x"829da433",
          8051 => x"70822b81",
          8052 => x"ffa41108",
          8053 => x"7033525c",
          8054 => x"56565673",
          8055 => x"762e8d38",
          8056 => x"8116701a",
          8057 => x"70335155",
          8058 => x"5673f538",
          8059 => x"82165473",
          8060 => x"7826a738",
          8061 => x"80557476",
          8062 => x"27913874",
          8063 => x"19547333",
          8064 => x"7a708105",
          8065 => x"5c348115",
          8066 => x"55ec39ba",
          8067 => x"7a708105",
          8068 => x"5c3474ff",
          8069 => x"2e098106",
          8070 => x"85389157",
          8071 => x"94396e18",
          8072 => x"81195954",
          8073 => x"73337a70",
          8074 => x"81055c34",
          8075 => x"7a7826ee",
          8076 => x"38807a34",
          8077 => x"768285ec",
          8078 => x"0c9e3d0d",
          8079 => x"04f73d0d",
          8080 => x"7b7d8d3d",
          8081 => x"fc055471",
          8082 => x"535755ec",
          8083 => x"ba3f8285",
          8084 => x"ec085382",
          8085 => x"85ec0882",
          8086 => x"fc389115",
          8087 => x"33537282",
          8088 => x"f4388c15",
          8089 => x"08547376",
          8090 => x"27923890",
          8091 => x"15337081",
          8092 => x"2a708106",
          8093 => x"51545772",
          8094 => x"83387356",
          8095 => x"94150854",
          8096 => x"80709417",
          8097 => x"0c587578",
          8098 => x"2e829938",
          8099 => x"798a1122",
          8100 => x"70892b59",
          8101 => x"51537378",
          8102 => x"2eb93876",
          8103 => x"52ff1651",
          8104 => x"fee0e73f",
          8105 => x"8285ec08",
          8106 => x"ff157854",
          8107 => x"70535553",
          8108 => x"fee0d73f",
          8109 => x"8285ec08",
          8110 => x"73269838",
          8111 => x"76098105",
          8112 => x"70750670",
          8113 => x"94180c77",
          8114 => x"71319818",
          8115 => x"08575851",
          8116 => x"53b13988",
          8117 => x"15085473",
          8118 => x"a6387352",
          8119 => x"7451cda0",
          8120 => x"3f8285ec",
          8121 => x"08548285",
          8122 => x"ec08812e",
          8123 => x"819a3882",
          8124 => x"85ec08ff",
          8125 => x"2e819b38",
          8126 => x"8285ec08",
          8127 => x"88160c73",
          8128 => x"98160c73",
          8129 => x"802e819c",
          8130 => x"38767627",
          8131 => x"80dc3875",
          8132 => x"77319416",
          8133 => x"08189417",
          8134 => x"0c901633",
          8135 => x"70812a70",
          8136 => x"81065155",
          8137 => x"5a567280",
          8138 => x"2e9a3873",
          8139 => x"527451cc",
          8140 => x"cf3f8285",
          8141 => x"ec085482",
          8142 => x"85ec0894",
          8143 => x"388285ec",
          8144 => x"0856a739",
          8145 => x"73527451",
          8146 => x"c6da3f82",
          8147 => x"85ec0854",
          8148 => x"73ff2ebe",
          8149 => x"38817427",
          8150 => x"af387953",
          8151 => x"73981408",
          8152 => x"27a63873",
          8153 => x"98160cff",
          8154 => x"a0399415",
          8155 => x"08169416",
          8156 => x"0c7583ff",
          8157 => x"06537280",
          8158 => x"2eaa3873",
          8159 => x"527951c5",
          8160 => x"f23f8285",
          8161 => x"ec089438",
          8162 => x"820b9116",
          8163 => x"34825380",
          8164 => x"c439810b",
          8165 => x"91163481",
          8166 => x"53bb3975",
          8167 => x"892a8285",
          8168 => x"ec080558",
          8169 => x"94150854",
          8170 => x"8c150874",
          8171 => x"27903873",
          8172 => x"8c160c90",
          8173 => x"153380c0",
          8174 => x"07537290",
          8175 => x"16347383",
          8176 => x"ff065372",
          8177 => x"802e8c38",
          8178 => x"779c1608",
          8179 => x"2e853877",
          8180 => x"9c160c80",
          8181 => x"53728285",
          8182 => x"ec0c8b3d",
          8183 => x"0d04f93d",
          8184 => x"0d795689",
          8185 => x"5475802e",
          8186 => x"818a3880",
          8187 => x"53893dfc",
          8188 => x"05528a3d",
          8189 => x"840551e1",
          8190 => x"dd3f8285",
          8191 => x"ec085582",
          8192 => x"85ec0880",
          8193 => x"ea387776",
          8194 => x"0c7a5275",
          8195 => x"51d8933f",
          8196 => x"8285ec08",
          8197 => x"558285ec",
          8198 => x"0880c338",
          8199 => x"ab163370",
          8200 => x"982b5557",
          8201 => x"807424a2",
          8202 => x"38861633",
          8203 => x"70842a70",
          8204 => x"81065155",
          8205 => x"5773802e",
          8206 => x"ad389c16",
          8207 => x"08527751",
          8208 => x"d3b83f82",
          8209 => x"85ec0888",
          8210 => x"170c7754",
          8211 => x"86142284",
          8212 => x"17237452",
          8213 => x"7551cec3",
          8214 => x"3f8285ec",
          8215 => x"08557484",
          8216 => x"2e098106",
          8217 => x"85388555",
          8218 => x"86397480",
          8219 => x"2e843880",
          8220 => x"760c7454",
          8221 => x"738285ec",
          8222 => x"0c893d0d",
          8223 => x"04fc3d0d",
          8224 => x"76873dfc",
          8225 => x"05537052",
          8226 => x"53e7fc3f",
          8227 => x"8285ec08",
          8228 => x"87388285",
          8229 => x"ec08730c",
          8230 => x"863d0d04",
          8231 => x"fb3d0d77",
          8232 => x"79893dfc",
          8233 => x"05547153",
          8234 => x"5654e7db",
          8235 => x"3f8285ec",
          8236 => x"08538285",
          8237 => x"ec0880e1",
          8238 => x"38749338",
          8239 => x"8285ec08",
          8240 => x"527351cd",
          8241 => x"d63f8285",
          8242 => x"ec085380",
          8243 => x"cc398285",
          8244 => x"ec085273",
          8245 => x"51d38a3f",
          8246 => x"8285ec08",
          8247 => x"538285ec",
          8248 => x"08842e09",
          8249 => x"81068538",
          8250 => x"80538739",
          8251 => x"8285ec08",
          8252 => x"a8387452",
          8253 => x"7351d591",
          8254 => x"3f725273",
          8255 => x"51cee73f",
          8256 => x"8285ec08",
          8257 => x"84327009",
          8258 => x"81057072",
          8259 => x"079f2c70",
          8260 => x"8285ec08",
          8261 => x"06515154",
          8262 => x"54728285",
          8263 => x"ec0c873d",
          8264 => x"0d04ee3d",
          8265 => x"0d655780",
          8266 => x"53893d70",
          8267 => x"53963d52",
          8268 => x"56dfa33f",
          8269 => x"8285ec08",
          8270 => x"558285ec",
          8271 => x"08b23864",
          8272 => x"527551d5",
          8273 => x"dd3f8285",
          8274 => x"ec085582",
          8275 => x"85ec08a0",
          8276 => x"380280cb",
          8277 => x"05337098",
          8278 => x"2b555873",
          8279 => x"80258538",
          8280 => x"86558d39",
          8281 => x"76802e88",
          8282 => x"38765275",
          8283 => x"51d49a3f",
          8284 => x"748285ec",
          8285 => x"0c943d0d",
          8286 => x"04f03d0d",
          8287 => x"6365555c",
          8288 => x"8053923d",
          8289 => x"ec055293",
          8290 => x"3d51deca",
          8291 => x"3f8285ec",
          8292 => x"085b8285",
          8293 => x"ec088287",
          8294 => x"387c740c",
          8295 => x"73089811",
          8296 => x"08fe1190",
          8297 => x"13085956",
          8298 => x"58557574",
          8299 => x"26913875",
          8300 => x"7c0c81eb",
          8301 => x"39815b81",
          8302 => x"d339825b",
          8303 => x"81ce3982",
          8304 => x"85ec0875",
          8305 => x"33555973",
          8306 => x"812e0981",
          8307 => x"0680c138",
          8308 => x"82755f57",
          8309 => x"7652923d",
          8310 => x"f00551c1",
          8311 => x"c73f8285",
          8312 => x"ec08ff2e",
          8313 => x"d0388285",
          8314 => x"ec08812e",
          8315 => x"cd388285",
          8316 => x"ec080981",
          8317 => x"05708285",
          8318 => x"ec080780",
          8319 => x"257a0581",
          8320 => x"197f5359",
          8321 => x"5a549814",
          8322 => x"087726c8",
          8323 => x"3880fd39",
          8324 => x"a4150882",
          8325 => x"85ec0857",
          8326 => x"58759838",
          8327 => x"77528118",
          8328 => x"7d5258ff",
          8329 => x"bed73f82",
          8330 => x"85ec085b",
          8331 => x"8285ec08",
          8332 => x"80da387c",
          8333 => x"70337712",
          8334 => x"ff1a5d52",
          8335 => x"56547482",
          8336 => x"2e098106",
          8337 => x"a038b414",
          8338 => x"51ffbb95",
          8339 => x"3f8285ec",
          8340 => x"0883ffff",
          8341 => x"06700981",
          8342 => x"05708025",
          8343 => x"1b821959",
          8344 => x"5b51549d",
          8345 => x"39b41451",
          8346 => x"ffbb8d3f",
          8347 => x"8285ec08",
          8348 => x"f00a0670",
          8349 => x"09810570",
          8350 => x"80251b84",
          8351 => x"19595b51",
          8352 => x"547583ff",
          8353 => x"067a5856",
          8354 => x"79ff8e38",
          8355 => x"787c0c7c",
          8356 => x"7990120c",
          8357 => x"84113381",
          8358 => x"07565474",
          8359 => x"8415347a",
          8360 => x"8285ec0c",
          8361 => x"923d0d04",
          8362 => x"f93d0d79",
          8363 => x"8a3dfc05",
          8364 => x"53705257",
          8365 => x"e3d13f82",
          8366 => x"85ec0856",
          8367 => x"8285ec08",
          8368 => x"81a83891",
          8369 => x"17335675",
          8370 => x"81a03890",
          8371 => x"17337081",
          8372 => x"2a708106",
          8373 => x"51555587",
          8374 => x"5573802e",
          8375 => x"818e3894",
          8376 => x"17085473",
          8377 => x"8c180827",
          8378 => x"81803873",
          8379 => x"9b388285",
          8380 => x"ec085388",
          8381 => x"17085276",
          8382 => x"51c3d93f",
          8383 => x"8285ec08",
          8384 => x"7488190c",
          8385 => x"5680c939",
          8386 => x"98170852",
          8387 => x"7651ffbf",
          8388 => x"933f8285",
          8389 => x"ec08ff2e",
          8390 => x"09810683",
          8391 => x"38815682",
          8392 => x"85ec0881",
          8393 => x"2e098106",
          8394 => x"85388256",
          8395 => x"a33975a0",
          8396 => x"38775482",
          8397 => x"85ec0898",
          8398 => x"15082794",
          8399 => x"38981708",
          8400 => x"538285ec",
          8401 => x"08527651",
          8402 => x"c38a3f82",
          8403 => x"85ec0856",
          8404 => x"9417088c",
          8405 => x"180c9017",
          8406 => x"3380c007",
          8407 => x"54739018",
          8408 => x"3475802e",
          8409 => x"85387591",
          8410 => x"18347555",
          8411 => x"748285ec",
          8412 => x"0c893d0d",
          8413 => x"04e23d0d",
          8414 => x"8253a03d",
          8415 => x"ffa40552",
          8416 => x"a13d51da",
          8417 => x"d13f8285",
          8418 => x"ec085582",
          8419 => x"85ec0881",
          8420 => x"f7387845",
          8421 => x"a13d0852",
          8422 => x"953d7052",
          8423 => x"58d1833f",
          8424 => x"8285ec08",
          8425 => x"558285ec",
          8426 => x"0881dd38",
          8427 => x"0280fb05",
          8428 => x"3370852a",
          8429 => x"70810651",
          8430 => x"55568655",
          8431 => x"7381c938",
          8432 => x"75982b54",
          8433 => x"80742481",
          8434 => x"bf380280",
          8435 => x"d6053370",
          8436 => x"81065854",
          8437 => x"87557681",
          8438 => x"af386b52",
          8439 => x"7851cc9a",
          8440 => x"3f8285ec",
          8441 => x"0874842a",
          8442 => x"70810651",
          8443 => x"55567380",
          8444 => x"2e80d438",
          8445 => x"78548285",
          8446 => x"ec089415",
          8447 => x"082e8188",
          8448 => x"38735a82",
          8449 => x"85ec085c",
          8450 => x"76528a3d",
          8451 => x"705254c7",
          8452 => x"8a3f8285",
          8453 => x"ec085582",
          8454 => x"85ec0880",
          8455 => x"eb388285",
          8456 => x"ec085273",
          8457 => x"51ccba3f",
          8458 => x"8285ec08",
          8459 => x"558285ec",
          8460 => x"08863887",
          8461 => x"5580d139",
          8462 => x"8285ec08",
          8463 => x"842e8838",
          8464 => x"8285ec08",
          8465 => x"80c23877",
          8466 => x"51ce973f",
          8467 => x"8285ec08",
          8468 => x"8285ec08",
          8469 => x"09810570",
          8470 => x"8285ec08",
          8471 => x"07802551",
          8472 => x"55557580",
          8473 => x"2e943873",
          8474 => x"802e8f38",
          8475 => x"80537552",
          8476 => x"7751c0e0",
          8477 => x"3f8285ec",
          8478 => x"0855748c",
          8479 => x"387851ff",
          8480 => x"bac23f82",
          8481 => x"85ec0855",
          8482 => x"748285ec",
          8483 => x"0ca03d0d",
          8484 => x"04e93d0d",
          8485 => x"8253993d",
          8486 => x"c005529a",
          8487 => x"3d51d8b6",
          8488 => x"3f8285ec",
          8489 => x"08548285",
          8490 => x"ec0882b0",
          8491 => x"38785e69",
          8492 => x"528e3d70",
          8493 => x"5258ceea",
          8494 => x"3f8285ec",
          8495 => x"08548285",
          8496 => x"ec088638",
          8497 => x"88548294",
          8498 => x"398285ec",
          8499 => x"08842e09",
          8500 => x"81068288",
          8501 => x"380280df",
          8502 => x"05337085",
          8503 => x"2a810651",
          8504 => x"55865474",
          8505 => x"81f63878",
          8506 => x"5a74528a",
          8507 => x"3d705257",
          8508 => x"c18e3f82",
          8509 => x"85ec0875",
          8510 => x"55568285",
          8511 => x"ec088338",
          8512 => x"87548285",
          8513 => x"ec08812e",
          8514 => x"09810683",
          8515 => x"38825482",
          8516 => x"85ec08ff",
          8517 => x"2e098106",
          8518 => x"86388154",
          8519 => x"81b43973",
          8520 => x"81b03882",
          8521 => x"85ec0852",
          8522 => x"7851c3f5",
          8523 => x"3f8285ec",
          8524 => x"08548285",
          8525 => x"ec08819a",
          8526 => x"388b53a0",
          8527 => x"52b41951",
          8528 => x"ffb6d03f",
          8529 => x"7854ae0b",
          8530 => x"b4153478",
          8531 => x"54900bbf",
          8532 => x"15348288",
          8533 => x"b20a5280",
          8534 => x"ca1951ff",
          8535 => x"b5e33f75",
          8536 => x"5378b411",
          8537 => x"5351c9cb",
          8538 => x"3fa05378",
          8539 => x"b4115380",
          8540 => x"d40551ff",
          8541 => x"b5fa3f78",
          8542 => x"54ae0b80",
          8543 => x"d515347f",
          8544 => x"537880d4",
          8545 => x"115351c9",
          8546 => x"aa3f7854",
          8547 => x"810b8315",
          8548 => x"347751ca",
          8549 => x"f73f8285",
          8550 => x"ec085482",
          8551 => x"85ec08b2",
          8552 => x"388288b2",
          8553 => x"0a526496",
          8554 => x"0551ffb5",
          8555 => x"943f7553",
          8556 => x"64527851",
          8557 => x"c8fd3f64",
          8558 => x"54900b8b",
          8559 => x"15347854",
          8560 => x"810b8315",
          8561 => x"347851ff",
          8562 => x"b7fa3f82",
          8563 => x"85ec0854",
          8564 => x"8b398053",
          8565 => x"75527651",
          8566 => x"ffbdf93f",
          8567 => x"738285ec",
          8568 => x"0c993d0d",
          8569 => x"04da3d0d",
          8570 => x"a93d8405",
          8571 => x"51d2d43f",
          8572 => x"8253a83d",
          8573 => x"ff840552",
          8574 => x"a93d51d5",
          8575 => x"d93f8285",
          8576 => x"ec085582",
          8577 => x"85ec0882",
          8578 => x"d338784d",
          8579 => x"a93d0852",
          8580 => x"9d3d7052",
          8581 => x"58cc8b3f",
          8582 => x"8285ec08",
          8583 => x"558285ec",
          8584 => x"0882b938",
          8585 => x"02819b05",
          8586 => x"3381a006",
          8587 => x"54865573",
          8588 => x"82aa38a0",
          8589 => x"53a43d08",
          8590 => x"52a83dff",
          8591 => x"880551ff",
          8592 => x"b4ae3fac",
          8593 => x"53775292",
          8594 => x"3d705254",
          8595 => x"ffb4a13f",
          8596 => x"aa3d0852",
          8597 => x"7351cbca",
          8598 => x"3f8285ec",
          8599 => x"08558285",
          8600 => x"ec089538",
          8601 => x"636f2e09",
          8602 => x"81068838",
          8603 => x"65a23d08",
          8604 => x"2e923888",
          8605 => x"5581e539",
          8606 => x"8285ec08",
          8607 => x"842e0981",
          8608 => x"0681b838",
          8609 => x"7351c984",
          8610 => x"3f8285ec",
          8611 => x"08558285",
          8612 => x"ec0881c8",
          8613 => x"38685693",
          8614 => x"53a83dff",
          8615 => x"9505528d",
          8616 => x"1651ffb3",
          8617 => x"cb3f02af",
          8618 => x"05338b17",
          8619 => x"348b1633",
          8620 => x"70842a70",
          8621 => x"81065155",
          8622 => x"55738938",
          8623 => x"74a00754",
          8624 => x"738b1734",
          8625 => x"7854810b",
          8626 => x"8315348b",
          8627 => x"16337084",
          8628 => x"2a708106",
          8629 => x"51555573",
          8630 => x"802e80e5",
          8631 => x"386e642e",
          8632 => x"80df3875",
          8633 => x"527851c6",
          8634 => x"913f8285",
          8635 => x"ec085278",
          8636 => x"51ffb6ff",
          8637 => x"3f825582",
          8638 => x"85ec0880",
          8639 => x"2e80dd38",
          8640 => x"8285ec08",
          8641 => x"527851ff",
          8642 => x"b4f33f82",
          8643 => x"85ec0879",
          8644 => x"80d41158",
          8645 => x"58558285",
          8646 => x"ec0880c0",
          8647 => x"38811633",
          8648 => x"5473ae2e",
          8649 => x"09810699",
          8650 => x"38635375",
          8651 => x"527651c6",
          8652 => x"823f7854",
          8653 => x"810b8315",
          8654 => x"34873982",
          8655 => x"85ec089c",
          8656 => x"387751c8",
          8657 => x"9d3f8285",
          8658 => x"ec085582",
          8659 => x"85ec088c",
          8660 => x"387851ff",
          8661 => x"b4ee3f82",
          8662 => x"85ec0855",
          8663 => x"748285ec",
          8664 => x"0ca83d0d",
          8665 => x"04ed3d0d",
          8666 => x"0280db05",
          8667 => x"33028405",
          8668 => x"80df0533",
          8669 => x"57578253",
          8670 => x"953dd005",
          8671 => x"52963d51",
          8672 => x"d2d43f82",
          8673 => x"85ec0855",
          8674 => x"8285ec08",
          8675 => x"80cf3878",
          8676 => x"5a655295",
          8677 => x"3dd40551",
          8678 => x"c9883f82",
          8679 => x"85ec0855",
          8680 => x"8285ec08",
          8681 => x"b8380280",
          8682 => x"cf053381",
          8683 => x"a0065486",
          8684 => x"5573aa38",
          8685 => x"75a70661",
          8686 => x"71098b12",
          8687 => x"3371067a",
          8688 => x"74060751",
          8689 => x"57555674",
          8690 => x"8b153478",
          8691 => x"54810b83",
          8692 => x"15347851",
          8693 => x"ffb3ed3f",
          8694 => x"8285ec08",
          8695 => x"55748285",
          8696 => x"ec0c953d",
          8697 => x"0d04ef3d",
          8698 => x"0d645682",
          8699 => x"53933dd0",
          8700 => x"0552943d",
          8701 => x"51d1df3f",
          8702 => x"8285ec08",
          8703 => x"558285ec",
          8704 => x"0880cb38",
          8705 => x"76586352",
          8706 => x"933dd405",
          8707 => x"51c8933f",
          8708 => x"8285ec08",
          8709 => x"558285ec",
          8710 => x"08b43802",
          8711 => x"80c70533",
          8712 => x"81a00654",
          8713 => x"865573a6",
          8714 => x"38841622",
          8715 => x"86172271",
          8716 => x"902b0753",
          8717 => x"54961f51",
          8718 => x"ffb0863f",
          8719 => x"7654810b",
          8720 => x"83153476",
          8721 => x"51ffb2fc",
          8722 => x"3f8285ec",
          8723 => x"08557482",
          8724 => x"85ec0c93",
          8725 => x"3d0d04ea",
          8726 => x"3d0d696b",
          8727 => x"5c5a8053",
          8728 => x"983dd005",
          8729 => x"52993d51",
          8730 => x"d0ec3f82",
          8731 => x"85ec0882",
          8732 => x"85ec0809",
          8733 => x"81057082",
          8734 => x"85ec0807",
          8735 => x"80255155",
          8736 => x"5779802e",
          8737 => x"81853881",
          8738 => x"70750655",
          8739 => x"5573802e",
          8740 => x"80f9387b",
          8741 => x"5d805f80",
          8742 => x"528d3d70",
          8743 => x"5254ffbd",
          8744 => x"fa3f8285",
          8745 => x"ec085782",
          8746 => x"85ec0880",
          8747 => x"d1387452",
          8748 => x"7351c3ad",
          8749 => x"3f8285ec",
          8750 => x"08578285",
          8751 => x"ec08bf38",
          8752 => x"8285ec08",
          8753 => x"8285ec08",
          8754 => x"655b5956",
          8755 => x"78188119",
          8756 => x"7b185659",
          8757 => x"55743374",
          8758 => x"34811656",
          8759 => x"8a7827ec",
          8760 => x"388b5675",
          8761 => x"1a548074",
          8762 => x"3475802e",
          8763 => x"9e38ff16",
          8764 => x"701b7033",
          8765 => x"51555673",
          8766 => x"a02ee838",
          8767 => x"8e397684",
          8768 => x"2e098106",
          8769 => x"8638807a",
          8770 => x"34805776",
          8771 => x"09810570",
          8772 => x"78078025",
          8773 => x"51547a80",
          8774 => x"2e80c138",
          8775 => x"73802ebc",
          8776 => x"387ba011",
          8777 => x"085351ff",
          8778 => x"b0d33f82",
          8779 => x"85ec0857",
          8780 => x"8285ec08",
          8781 => x"a7387b70",
          8782 => x"33555580",
          8783 => x"c3567383",
          8784 => x"2e8b3880",
          8785 => x"e4567384",
          8786 => x"2e8338a7",
          8787 => x"567515b4",
          8788 => x"0551ffad",
          8789 => x"a33f8285",
          8790 => x"ec087b0c",
          8791 => x"768285ec",
          8792 => x"0c983d0d",
          8793 => x"04e63d0d",
          8794 => x"82539c3d",
          8795 => x"ffb80552",
          8796 => x"9d3d51ce",
          8797 => x"e13f8285",
          8798 => x"ec088285",
          8799 => x"ec085654",
          8800 => x"8285ec08",
          8801 => x"8398388b",
          8802 => x"53a0528b",
          8803 => x"3d705259",
          8804 => x"ffae803f",
          8805 => x"736d7033",
          8806 => x"7081ff06",
          8807 => x"52575557",
          8808 => x"9f742781",
          8809 => x"bc387858",
          8810 => x"7481ff06",
          8811 => x"6d81054e",
          8812 => x"705255ff",
          8813 => x"aec93f82",
          8814 => x"85ec0880",
          8815 => x"2ea5386c",
          8816 => x"70337053",
          8817 => x"5754ffae",
          8818 => x"bd3f8285",
          8819 => x"ec08802e",
          8820 => x"8d387488",
          8821 => x"2b76076d",
          8822 => x"81054e55",
          8823 => x"86398285",
          8824 => x"ec0855ff",
          8825 => x"9f157083",
          8826 => x"ffff0651",
          8827 => x"54739926",
          8828 => x"8a38e015",
          8829 => x"7083ffff",
          8830 => x"06565480",
          8831 => x"ff752787",
          8832 => x"3881feb4",
          8833 => x"15335574",
          8834 => x"802ea338",
          8835 => x"74528280",
          8836 => x"b451ffad",
          8837 => x"c93f8285",
          8838 => x"ec089338",
          8839 => x"81ff7527",
          8840 => x"88387689",
          8841 => x"2688388b",
          8842 => x"398a7727",
          8843 => x"86388655",
          8844 => x"81ec3981",
          8845 => x"ff75278f",
          8846 => x"3874882a",
          8847 => x"54737870",
          8848 => x"81055a34",
          8849 => x"81175774",
          8850 => x"78708105",
          8851 => x"5a348117",
          8852 => x"6d703370",
          8853 => x"81ff0652",
          8854 => x"57555773",
          8855 => x"9f26fec8",
          8856 => x"388b3d33",
          8857 => x"54865573",
          8858 => x"81e52e81",
          8859 => x"b1387680",
          8860 => x"2e993802",
          8861 => x"a7055576",
          8862 => x"15703351",
          8863 => x"5473a02e",
          8864 => x"09810687",
          8865 => x"38ff1757",
          8866 => x"76ed3879",
          8867 => x"41804380",
          8868 => x"52913d70",
          8869 => x"5255ffba",
          8870 => x"823f8285",
          8871 => x"ec085482",
          8872 => x"85ec0880",
          8873 => x"f7388152",
          8874 => x"7451ffbf",
          8875 => x"b43f8285",
          8876 => x"ec085482",
          8877 => x"85ec088d",
          8878 => x"387680c4",
          8879 => x"386754e5",
          8880 => x"743480c6",
          8881 => x"398285ec",
          8882 => x"08842e09",
          8883 => x"810680cc",
          8884 => x"38805476",
          8885 => x"742e80c4",
          8886 => x"38815274",
          8887 => x"51ffbcff",
          8888 => x"3f8285ec",
          8889 => x"08548285",
          8890 => x"ec08b138",
          8891 => x"a0538285",
          8892 => x"ec085267",
          8893 => x"51ffab9b",
          8894 => x"3f675488",
          8895 => x"0b8b1534",
          8896 => x"8b537852",
          8897 => x"6751ffaa",
          8898 => x"e73f7954",
          8899 => x"810b8315",
          8900 => x"347951ff",
          8901 => x"adae3f82",
          8902 => x"85ec0854",
          8903 => x"73557482",
          8904 => x"85ec0c9c",
          8905 => x"3d0d04f2",
          8906 => x"3d0d6062",
          8907 => x"02880580",
          8908 => x"cb053393",
          8909 => x"3dfc0555",
          8910 => x"7254405e",
          8911 => x"5ad2c83f",
          8912 => x"8285ec08",
          8913 => x"588285ec",
          8914 => x"0882bf38",
          8915 => x"911a3358",
          8916 => x"7782b738",
          8917 => x"7c802e97",
          8918 => x"388c1a08",
          8919 => x"59789038",
          8920 => x"901a3370",
          8921 => x"812a7081",
          8922 => x"06515555",
          8923 => x"73903887",
          8924 => x"54829939",
          8925 => x"82588292",
          8926 => x"39815882",
          8927 => x"8d397e8a",
          8928 => x"11227089",
          8929 => x"2b70557f",
          8930 => x"54565656",
          8931 => x"fec6fb3f",
          8932 => x"ff147d06",
          8933 => x"70098105",
          8934 => x"7072079f",
          8935 => x"2a8285ec",
          8936 => x"08058c19",
          8937 => x"087c405a",
          8938 => x"5d555581",
          8939 => x"77278838",
          8940 => x"98160877",
          8941 => x"26833882",
          8942 => x"57767756",
          8943 => x"59805674",
          8944 => x"527951ff",
          8945 => x"adde3f81",
          8946 => x"157f5555",
          8947 => x"98140875",
          8948 => x"26833882",
          8949 => x"558285ec",
          8950 => x"08812eff",
          8951 => x"97388285",
          8952 => x"ec08ff2e",
          8953 => x"ff933882",
          8954 => x"85ec088e",
          8955 => x"38811656",
          8956 => x"757b2e09",
          8957 => x"81068738",
          8958 => x"93397459",
          8959 => x"80567477",
          8960 => x"2e098106",
          8961 => x"ffb93887",
          8962 => x"5880ff39",
          8963 => x"7d802eba",
          8964 => x"38787b55",
          8965 => x"557a802e",
          8966 => x"b4388115",
          8967 => x"5673812e",
          8968 => x"09810683",
          8969 => x"38ff5675",
          8970 => x"5374527e",
          8971 => x"51ffaeed",
          8972 => x"3f8285ec",
          8973 => x"08588285",
          8974 => x"ec0880ce",
          8975 => x"38748116",
          8976 => x"ff165656",
          8977 => x"5c73d338",
          8978 => x"8439ff19",
          8979 => x"5c7e7c8c",
          8980 => x"120c557d",
          8981 => x"802eb338",
          8982 => x"78881b0c",
          8983 => x"7c8c1b0c",
          8984 => x"901a3380",
          8985 => x"c0075473",
          8986 => x"901b3498",
          8987 => x"1508fe05",
          8988 => x"90160857",
          8989 => x"54757426",
          8990 => x"9138757b",
          8991 => x"3190160c",
          8992 => x"84153381",
          8993 => x"07547384",
          8994 => x"16347754",
          8995 => x"738285ec",
          8996 => x"0c903d0d",
          8997 => x"04e93d0d",
          8998 => x"6b6d0288",
          8999 => x"0580eb05",
          9000 => x"339d3d54",
          9001 => x"5a5c59c5",
          9002 => x"9a3f8b56",
          9003 => x"800b8285",
          9004 => x"ec08248c",
          9005 => x"82388285",
          9006 => x"ec08822b",
          9007 => x"829d9011",
          9008 => x"08515574",
          9009 => x"802e8438",
          9010 => x"80753482",
          9011 => x"85ec0881",
          9012 => x"ff065f81",
          9013 => x"527e51ff",
          9014 => x"a08f3f82",
          9015 => x"85ec0881",
          9016 => x"ff067081",
          9017 => x"06565783",
          9018 => x"56748bcb",
          9019 => x"3876822a",
          9020 => x"70810651",
          9021 => x"558a5674",
          9022 => x"8bbd3899",
          9023 => x"3dfc0553",
          9024 => x"83527e51",
          9025 => x"ffa4af3f",
          9026 => x"8285ec08",
          9027 => x"99386755",
          9028 => x"74802e92",
          9029 => x"38748280",
          9030 => x"80268b38",
          9031 => x"ff157506",
          9032 => x"5574802e",
          9033 => x"83388148",
          9034 => x"78802e87",
          9035 => x"38848079",
          9036 => x"26923878",
          9037 => x"81800a26",
          9038 => x"8b38ff19",
          9039 => x"79065574",
          9040 => x"802e8638",
          9041 => x"93568aef",
          9042 => x"3978892a",
          9043 => x"6e892a70",
          9044 => x"892b7759",
          9045 => x"4843597a",
          9046 => x"83388156",
          9047 => x"61098105",
          9048 => x"70802577",
          9049 => x"07515591",
          9050 => x"56748acb",
          9051 => x"38993df8",
          9052 => x"05538152",
          9053 => x"7e51ffa3",
          9054 => x"bd3f8156",
          9055 => x"8285ec08",
          9056 => x"8ab53877",
          9057 => x"832a7077",
          9058 => x"068285ec",
          9059 => x"08435645",
          9060 => x"748338bf",
          9061 => x"4166558e",
          9062 => x"56607526",
          9063 => x"8a993874",
          9064 => x"61317048",
          9065 => x"5580ff75",
          9066 => x"278a8c38",
          9067 => x"93567881",
          9068 => x"80268a83",
          9069 => x"3877812a",
          9070 => x"70810656",
          9071 => x"4374802e",
          9072 => x"95387787",
          9073 => x"06557482",
          9074 => x"2e839438",
          9075 => x"77810655",
          9076 => x"74802e83",
          9077 => x"8a387781",
          9078 => x"06559356",
          9079 => x"825e7480",
          9080 => x"2e89d438",
          9081 => x"785a7d83",
          9082 => x"2e098106",
          9083 => x"80e03878",
          9084 => x"ae386691",
          9085 => x"2a57810b",
          9086 => x"8280d822",
          9087 => x"565a7480",
          9088 => x"2e9d3874",
          9089 => x"77269838",
          9090 => x"8280d856",
          9091 => x"79108217",
          9092 => x"70225757",
          9093 => x"5a74802e",
          9094 => x"86387675",
          9095 => x"27ee3879",
          9096 => x"526651fe",
          9097 => x"c1e43f82",
          9098 => x"85ec0882",
          9099 => x"2b848711",
          9100 => x"892a5e55",
          9101 => x"a05c800b",
          9102 => x"8285ec08",
          9103 => x"fc808a05",
          9104 => x"5644fdff",
          9105 => x"f00a7527",
          9106 => x"80f23888",
          9107 => x"dd3978ae",
          9108 => x"38668c2a",
          9109 => x"57810b82",
          9110 => x"80c82256",
          9111 => x"5a74802e",
          9112 => x"9d387477",
          9113 => x"26983882",
          9114 => x"80c85679",
          9115 => x"10821770",
          9116 => x"2257575a",
          9117 => x"74802e86",
          9118 => x"38767527",
          9119 => x"ee387952",
          9120 => x"6651fec1",
          9121 => x"853f8285",
          9122 => x"ec088285",
          9123 => x"ec080584",
          9124 => x"05578285",
          9125 => x"ec089ff5",
          9126 => x"26983881",
          9127 => x"0b8285ec",
          9128 => x"08712b82",
          9129 => x"85ec0811",
          9130 => x"1270732a",
          9131 => x"83055a51",
          9132 => x"565e83ff",
          9133 => x"17892a5d",
          9134 => x"815ca044",
          9135 => x"601c7d11",
          9136 => x"65056970",
          9137 => x"12ff0571",
          9138 => x"09810570",
          9139 => x"72067431",
          9140 => x"5c525957",
          9141 => x"59407d83",
          9142 => x"2e098106",
          9143 => x"8938761c",
          9144 => x"6018415c",
          9145 => x"8439761d",
          9146 => x"5d79842b",
          9147 => x"70196231",
          9148 => x"68585155",
          9149 => x"74762687",
          9150 => x"b138757c",
          9151 => x"317d317a",
          9152 => x"53706531",
          9153 => x"5255fec0",
          9154 => x"813f8285",
          9155 => x"ec08587d",
          9156 => x"832e0981",
          9157 => x"069b3882",
          9158 => x"85ec0883",
          9159 => x"fff52680",
          9160 => x"dd387887",
          9161 => x"85387981",
          9162 => x"2a5978fd",
          9163 => x"b73886fa",
          9164 => x"397d822e",
          9165 => x"09810680",
          9166 => x"c53883ff",
          9167 => x"f50b8285",
          9168 => x"ec0827a0",
          9169 => x"38788f38",
          9170 => x"791a5574",
          9171 => x"80c02686",
          9172 => x"387459fd",
          9173 => x"8f396281",
          9174 => x"06557480",
          9175 => x"2e8f3883",
          9176 => x"5efd8139",
          9177 => x"8285ec08",
          9178 => x"9ff52692",
          9179 => x"387886ba",
          9180 => x"38791a59",
          9181 => x"81807927",
          9182 => x"fcea3886",
          9183 => x"ad398055",
          9184 => x"7d812e09",
          9185 => x"81068338",
          9186 => x"7d559ff5",
          9187 => x"78278b38",
          9188 => x"74810655",
          9189 => x"8e567486",
          9190 => x"9e388480",
          9191 => x"5380527a",
          9192 => x"51ffa1ef",
          9193 => x"3f8b5381",
          9194 => x"fef0527a",
          9195 => x"51ffa1c0",
          9196 => x"3f848052",
          9197 => x"8b1b51ff",
          9198 => x"a0e93f79",
          9199 => x"8d1c347b",
          9200 => x"83ffff06",
          9201 => x"528e1b51",
          9202 => x"ffa0d83f",
          9203 => x"810b901c",
          9204 => x"347d8332",
          9205 => x"70098105",
          9206 => x"70962a84",
          9207 => x"80065451",
          9208 => x"55911b51",
          9209 => x"ffa0bc3f",
          9210 => x"66557483",
          9211 => x"ffff2690",
          9212 => x"387483ff",
          9213 => x"ff065293",
          9214 => x"1b51ffa0",
          9215 => x"a63f8a39",
          9216 => x"7452a01b",
          9217 => x"51ffa0b9",
          9218 => x"3ff80b95",
          9219 => x"1c34bf52",
          9220 => x"981b51ff",
          9221 => x"a08d3f81",
          9222 => x"ff529a1b",
          9223 => x"51ffa083",
          9224 => x"3f60529c",
          9225 => x"1b51ffa0",
          9226 => x"983f7d83",
          9227 => x"2e098106",
          9228 => x"80cb3882",
          9229 => x"88b20a52",
          9230 => x"80c31b51",
          9231 => x"ffa0823f",
          9232 => x"7c52a41b",
          9233 => x"51ff9ff9",
          9234 => x"3f8252ac",
          9235 => x"1b51ff9f",
          9236 => x"f03f8152",
          9237 => x"b01b51ff",
          9238 => x"9fc93f86",
          9239 => x"52b21b51",
          9240 => x"ff9fc03f",
          9241 => x"ff800b80",
          9242 => x"c01c34a9",
          9243 => x"0b80c21c",
          9244 => x"34935381",
          9245 => x"fefc5280",
          9246 => x"c71b51ae",
          9247 => x"398288b2",
          9248 => x"0a52a71b",
          9249 => x"51ff9fb9",
          9250 => x"3f7c83ff",
          9251 => x"ff065296",
          9252 => x"1b51ff9f",
          9253 => x"8e3fff80",
          9254 => x"0ba41c34",
          9255 => x"a90ba61c",
          9256 => x"34935381",
          9257 => x"ff9052ab",
          9258 => x"1b51ff9f",
          9259 => x"c33f82d4",
          9260 => x"d55283fe",
          9261 => x"1b705259",
          9262 => x"ff9ee83f",
          9263 => x"81546053",
          9264 => x"7a527e51",
          9265 => x"ff9b8b3f",
          9266 => x"81568285",
          9267 => x"ec0883e7",
          9268 => x"387d832e",
          9269 => x"09810680",
          9270 => x"ee387554",
          9271 => x"60860553",
          9272 => x"7a527e51",
          9273 => x"ff9aeb3f",
          9274 => x"84805380",
          9275 => x"527a51ff",
          9276 => x"9fa13f84",
          9277 => x"8b85a4d2",
          9278 => x"527a51ff",
          9279 => x"9ec33f86",
          9280 => x"8a85e4f2",
          9281 => x"5283e41b",
          9282 => x"51ff9eb5",
          9283 => x"3fff1852",
          9284 => x"83e81b51",
          9285 => x"ff9eaa3f",
          9286 => x"825283ec",
          9287 => x"1b51ff9e",
          9288 => x"a03f82d4",
          9289 => x"d5527851",
          9290 => x"ff9df83f",
          9291 => x"75546087",
          9292 => x"05537a52",
          9293 => x"7e51ff9a",
          9294 => x"993f7554",
          9295 => x"6016537a",
          9296 => x"527e51ff",
          9297 => x"9a8c3f65",
          9298 => x"5380527a",
          9299 => x"51ff9ec3",
          9300 => x"3f7f5680",
          9301 => x"587d832e",
          9302 => x"0981069a",
          9303 => x"38f8527a",
          9304 => x"51ff9ddd",
          9305 => x"3fff5284",
          9306 => x"1b51ff9d",
          9307 => x"d43ff00a",
          9308 => x"52881b51",
          9309 => x"913987ff",
          9310 => x"fff8557d",
          9311 => x"812e8338",
          9312 => x"f8557452",
          9313 => x"7a51ff9d",
          9314 => x"b83f7c55",
          9315 => x"61577462",
          9316 => x"26833874",
          9317 => x"57765475",
          9318 => x"537a527e",
          9319 => x"51ff99b2",
          9320 => x"3f8285ec",
          9321 => x"08828738",
          9322 => x"84805382",
          9323 => x"85ec0852",
          9324 => x"7a51ff9d",
          9325 => x"de3f7616",
          9326 => x"75783156",
          9327 => x"5674cd38",
          9328 => x"81185877",
          9329 => x"802eff8d",
          9330 => x"3879557d",
          9331 => x"832e8338",
          9332 => x"63556157",
          9333 => x"74622683",
          9334 => x"38745776",
          9335 => x"5475537a",
          9336 => x"527e51ff",
          9337 => x"98ec3f82",
          9338 => x"85ec0881",
          9339 => x"c1387616",
          9340 => x"75783156",
          9341 => x"5674db38",
          9342 => x"8c567d83",
          9343 => x"2e933886",
          9344 => x"566683ff",
          9345 => x"ff268a38",
          9346 => x"84567d82",
          9347 => x"2e833881",
          9348 => x"56648106",
          9349 => x"587780fe",
          9350 => x"38848053",
          9351 => x"77527a51",
          9352 => x"ff9cf03f",
          9353 => x"82d4d552",
          9354 => x"7851ff9b",
          9355 => x"f63f83be",
          9356 => x"1b557775",
          9357 => x"34810b81",
          9358 => x"1634810b",
          9359 => x"82163477",
          9360 => x"83163475",
          9361 => x"84163460",
          9362 => x"67055680",
          9363 => x"fdc15275",
          9364 => x"51feb9b6",
          9365 => x"3ffe0b85",
          9366 => x"16348285",
          9367 => x"ec08822a",
          9368 => x"bf075675",
          9369 => x"86163482",
          9370 => x"85ec0887",
          9371 => x"16346052",
          9372 => x"83c61b51",
          9373 => x"ff9bca3f",
          9374 => x"665283ca",
          9375 => x"1b51ff9b",
          9376 => x"c03f8154",
          9377 => x"77537a52",
          9378 => x"7e51ff97",
          9379 => x"c53f8156",
          9380 => x"8285ec08",
          9381 => x"a2388053",
          9382 => x"80527e51",
          9383 => x"ff99973f",
          9384 => x"81568285",
          9385 => x"ec089038",
          9386 => x"89398e56",
          9387 => x"8a398156",
          9388 => x"86398285",
          9389 => x"ec085675",
          9390 => x"8285ec0c",
          9391 => x"993d0d04",
          9392 => x"f53d0d7d",
          9393 => x"605b5980",
          9394 => x"7960ff05",
          9395 => x"5a575776",
          9396 => x"7825b438",
          9397 => x"8d3df811",
          9398 => x"55558153",
          9399 => x"fc155279",
          9400 => x"51c9c03f",
          9401 => x"7a812e09",
          9402 => x"81069c38",
          9403 => x"8c3d3355",
          9404 => x"748d2edb",
          9405 => x"38747670",
          9406 => x"81055834",
          9407 => x"81175774",
          9408 => x"8a2e0981",
          9409 => x"06c93880",
          9410 => x"76347855",
          9411 => x"76833876",
          9412 => x"55748285",
          9413 => x"ec0c8d3d",
          9414 => x"0d04f73d",
          9415 => x"0d7b0284",
          9416 => x"05b30533",
          9417 => x"5957778a",
          9418 => x"2e098106",
          9419 => x"87388d52",
          9420 => x"7651e73f",
          9421 => x"84170856",
          9422 => x"80762480",
          9423 => x"c2388817",
          9424 => x"0877178c",
          9425 => x"05565977",
          9426 => x"75348116",
          9427 => x"56bb7625",
          9428 => x"a5388b3d",
          9429 => x"fc055475",
          9430 => x"538c1752",
          9431 => x"760851cb",
          9432 => x"bf3f7976",
          9433 => x"32700981",
          9434 => x"05707207",
          9435 => x"9f2a7009",
          9436 => x"81055351",
          9437 => x"56567584",
          9438 => x"180c8119",
          9439 => x"88180c8b",
          9440 => x"3d0d04f9",
          9441 => x"3d0d7984",
          9442 => x"11085656",
          9443 => x"807524a7",
          9444 => x"38893dfc",
          9445 => x"05547453",
          9446 => x"8c165275",
          9447 => x"0851cb80",
          9448 => x"3f8285ec",
          9449 => x"08913884",
          9450 => x"1608782e",
          9451 => x"09810687",
          9452 => x"38881608",
          9453 => x"558339ff",
          9454 => x"55748285",
          9455 => x"ec0c893d",
          9456 => x"0d04fd3d",
          9457 => x"0d755480",
          9458 => x"cc538052",
          9459 => x"7351ff99",
          9460 => x"c23f7674",
          9461 => x"0c853d0d",
          9462 => x"04ea3d0d",
          9463 => x"0280e305",
          9464 => x"336a5386",
          9465 => x"3d705354",
          9466 => x"54d83f73",
          9467 => x"527251fe",
          9468 => x"a93f7251",
          9469 => x"ff8d3f98",
          9470 => x"3d0d0400",
          9471 => x"00ffffff",
          9472 => x"ff00ffff",
          9473 => x"ffff00ff",
          9474 => x"ffffff00",
          9475 => x"0000118e",
          9476 => x"00001112",
          9477 => x"00001119",
          9478 => x"00001120",
          9479 => x"00001127",
          9480 => x"0000112e",
          9481 => x"00001135",
          9482 => x"0000113c",
          9483 => x"00001143",
          9484 => x"0000114a",
          9485 => x"00001151",
          9486 => x"00001158",
          9487 => x"0000115e",
          9488 => x"00001164",
          9489 => x"0000116a",
          9490 => x"00001170",
          9491 => x"00001176",
          9492 => x"0000117c",
          9493 => x"00001182",
          9494 => x"00001188",
          9495 => x"000026ce",
          9496 => x"000026d4",
          9497 => x"000026da",
          9498 => x"000026e0",
          9499 => x"000026e6",
          9500 => x"000032e6",
          9501 => x"000033d0",
          9502 => x"000034bd",
          9503 => x"000036eb",
          9504 => x"000033b8",
          9505 => x"000031c3",
          9506 => x"00003567",
          9507 => x"000036c2",
          9508 => x"000035a4",
          9509 => x"0000363b",
          9510 => x"000035c0",
          9511 => x"0000346d",
          9512 => x"000031c3",
          9513 => x"000034bd",
          9514 => x"000034e0",
          9515 => x"00003567",
          9516 => x"000031c3",
          9517 => x"000031c3",
          9518 => x"000035c0",
          9519 => x"0000363b",
          9520 => x"000036c2",
          9521 => x"000036eb",
          9522 => x"64696e69",
          9523 => x"74000000",
          9524 => x"64696f63",
          9525 => x"746c0000",
          9526 => x"66696e69",
          9527 => x"74000000",
          9528 => x"666c6f61",
          9529 => x"64000000",
          9530 => x"66657865",
          9531 => x"63000000",
          9532 => x"6d636c65",
          9533 => x"61720000",
          9534 => x"6d636f70",
          9535 => x"79000000",
          9536 => x"6d646966",
          9537 => x"66000000",
          9538 => x"6d64756d",
          9539 => x"70000000",
          9540 => x"6d656200",
          9541 => x"6d656800",
          9542 => x"6d657700",
          9543 => x"68696400",
          9544 => x"68696500",
          9545 => x"68666400",
          9546 => x"68666500",
          9547 => x"63616c6c",
          9548 => x"00000000",
          9549 => x"6a6d7000",
          9550 => x"72657374",
          9551 => x"61727400",
          9552 => x"72657365",
          9553 => x"74000000",
          9554 => x"696e666f",
          9555 => x"00000000",
          9556 => x"74657374",
          9557 => x"00000000",
          9558 => x"74626173",
          9559 => x"69630000",
          9560 => x"6d626173",
          9561 => x"69630000",
          9562 => x"6b696c6f",
          9563 => x"00000000",
          9564 => x"65640000",
          9565 => x"4469736b",
          9566 => x"20457272",
          9567 => x"6f720a00",
          9568 => x"496e7465",
          9569 => x"726e616c",
          9570 => x"20657272",
          9571 => x"6f722e0a",
          9572 => x"00000000",
          9573 => x"4469736b",
          9574 => x"206e6f74",
          9575 => x"20726561",
          9576 => x"64792e0a",
          9577 => x"00000000",
          9578 => x"4e6f2066",
          9579 => x"696c6520",
          9580 => x"666f756e",
          9581 => x"642e0a00",
          9582 => x"4e6f2070",
          9583 => x"61746820",
          9584 => x"666f756e",
          9585 => x"642e0a00",
          9586 => x"496e7661",
          9587 => x"6c696420",
          9588 => x"66696c65",
          9589 => x"6e616d65",
          9590 => x"2e0a0000",
          9591 => x"41636365",
          9592 => x"73732064",
          9593 => x"656e6965",
          9594 => x"642e0a00",
          9595 => x"46696c65",
          9596 => x"20616c72",
          9597 => x"65616479",
          9598 => x"20657869",
          9599 => x"7374732e",
          9600 => x"0a000000",
          9601 => x"46696c65",
          9602 => x"2068616e",
          9603 => x"646c6520",
          9604 => x"696e7661",
          9605 => x"6c69642e",
          9606 => x"0a000000",
          9607 => x"53442069",
          9608 => x"73207772",
          9609 => x"69746520",
          9610 => x"70726f74",
          9611 => x"65637465",
          9612 => x"642e0a00",
          9613 => x"44726976",
          9614 => x"65206e75",
          9615 => x"6d626572",
          9616 => x"20697320",
          9617 => x"696e7661",
          9618 => x"6c69642e",
          9619 => x"0a000000",
          9620 => x"4469736b",
          9621 => x"206e6f74",
          9622 => x"20656e61",
          9623 => x"626c6564",
          9624 => x"2e0a0000",
          9625 => x"4e6f2063",
          9626 => x"6f6d7061",
          9627 => x"7469626c",
          9628 => x"65206669",
          9629 => x"6c657379",
          9630 => x"7374656d",
          9631 => x"20666f75",
          9632 => x"6e64206f",
          9633 => x"6e206469",
          9634 => x"736b2e0a",
          9635 => x"00000000",
          9636 => x"466f726d",
          9637 => x"61742061",
          9638 => x"626f7274",
          9639 => x"65642e0a",
          9640 => x"00000000",
          9641 => x"54696d65",
          9642 => x"6f75742c",
          9643 => x"206f7065",
          9644 => x"72617469",
          9645 => x"6f6e2063",
          9646 => x"616e6365",
          9647 => x"6c6c6564",
          9648 => x"2e0a0000",
          9649 => x"46696c65",
          9650 => x"20697320",
          9651 => x"6c6f636b",
          9652 => x"65642e0a",
          9653 => x"00000000",
          9654 => x"496e7375",
          9655 => x"66666963",
          9656 => x"69656e74",
          9657 => x"206d656d",
          9658 => x"6f72792e",
          9659 => x"0a000000",
          9660 => x"546f6f20",
          9661 => x"6d616e79",
          9662 => x"206f7065",
          9663 => x"6e206669",
          9664 => x"6c65732e",
          9665 => x"0a000000",
          9666 => x"50617261",
          9667 => x"6d657465",
          9668 => x"72732069",
          9669 => x"6e636f72",
          9670 => x"72656374",
          9671 => x"2e0a0000",
          9672 => x"53756363",
          9673 => x"6573732e",
          9674 => x"0a000000",
          9675 => x"556e6b6e",
          9676 => x"6f776e20",
          9677 => x"6572726f",
          9678 => x"722e0a00",
          9679 => x"0a256c75",
          9680 => x"20627974",
          9681 => x"65732025",
          9682 => x"73206174",
          9683 => x"20256c75",
          9684 => x"20627974",
          9685 => x"65732f73",
          9686 => x"65632e0a",
          9687 => x"00000000",
          9688 => x"72656164",
          9689 => x"00000000",
          9690 => x"25303858",
          9691 => x"00000000",
          9692 => x"3a202000",
          9693 => x"25303458",
          9694 => x"00000000",
          9695 => x"20202020",
          9696 => x"20202020",
          9697 => x"00000000",
          9698 => x"25303258",
          9699 => x"00000000",
          9700 => x"20200000",
          9701 => x"207c0000",
          9702 => x"7c0d0a00",
          9703 => x"7a4f5300",
          9704 => x"0a2a2a20",
          9705 => x"25732028",
          9706 => x"00000000",
          9707 => x"30322f30",
          9708 => x"352f3230",
          9709 => x"32300000",
          9710 => x"76312e30",
          9711 => x"32000000",
          9712 => x"205a5055",
          9713 => x"2c207265",
          9714 => x"76202530",
          9715 => x"32782920",
          9716 => x"25732025",
          9717 => x"73202a2a",
          9718 => x"0a0a0000",
          9719 => x"5a505520",
          9720 => x"496e7465",
          9721 => x"72727570",
          9722 => x"74204861",
          9723 => x"6e646c65",
          9724 => x"720a0000",
          9725 => x"54696d65",
          9726 => x"7220696e",
          9727 => x"74657272",
          9728 => x"7570740a",
          9729 => x"00000000",
          9730 => x"50533220",
          9731 => x"696e7465",
          9732 => x"72727570",
          9733 => x"740a0000",
          9734 => x"494f4354",
          9735 => x"4c205244",
          9736 => x"20696e74",
          9737 => x"65727275",
          9738 => x"70740a00",
          9739 => x"494f4354",
          9740 => x"4c205752",
          9741 => x"20696e74",
          9742 => x"65727275",
          9743 => x"70740a00",
          9744 => x"55415254",
          9745 => x"30205258",
          9746 => x"20696e74",
          9747 => x"65727275",
          9748 => x"70740a00",
          9749 => x"55415254",
          9750 => x"30205458",
          9751 => x"20696e74",
          9752 => x"65727275",
          9753 => x"70740a00",
          9754 => x"55415254",
          9755 => x"31205258",
          9756 => x"20696e74",
          9757 => x"65727275",
          9758 => x"70740a00",
          9759 => x"55415254",
          9760 => x"31205458",
          9761 => x"20696e74",
          9762 => x"65727275",
          9763 => x"70740a00",
          9764 => x"53657474",
          9765 => x"696e6720",
          9766 => x"75702074",
          9767 => x"696d6572",
          9768 => x"2e2e2e0a",
          9769 => x"00000000",
          9770 => x"456e6162",
          9771 => x"6c696e67",
          9772 => x"2074696d",
          9773 => x"65722e2e",
          9774 => x"2e0a0000",
          9775 => x"6175746f",
          9776 => x"65786563",
          9777 => x"2e626174",
          9778 => x"00000000",
          9779 => x"7a4f532e",
          9780 => x"68737400",
          9781 => x"303a0000",
          9782 => x"4661696c",
          9783 => x"65642074",
          9784 => x"6f20696e",
          9785 => x"69746961",
          9786 => x"6c697365",
          9787 => x"20736420",
          9788 => x"63617264",
          9789 => x"20302c20",
          9790 => x"706c6561",
          9791 => x"73652069",
          9792 => x"6e697420",
          9793 => x"6d616e75",
          9794 => x"616c6c79",
          9795 => x"2e0a0000",
          9796 => x"2a200000",
          9797 => x"436c6561",
          9798 => x"72696e67",
          9799 => x"2e2e2e2e",
          9800 => x"00000000",
          9801 => x"436f7079",
          9802 => x"696e672e",
          9803 => x"2e2e0000",
          9804 => x"436f6d70",
          9805 => x"6172696e",
          9806 => x"672e2e2e",
          9807 => x"00000000",
          9808 => x"2530386c",
          9809 => x"78282530",
          9810 => x"3878292d",
          9811 => x"3e253038",
          9812 => x"6c782825",
          9813 => x"30387829",
          9814 => x"0a000000",
          9815 => x"44756d70",
          9816 => x"204d656d",
          9817 => x"6f72790a",
          9818 => x"00000000",
          9819 => x"0a436f6d",
          9820 => x"706c6574",
          9821 => x"652e0a00",
          9822 => x"25303858",
          9823 => x"20253032",
          9824 => x"582d0000",
          9825 => x"3f3f3f0a",
          9826 => x"00000000",
          9827 => x"25303858",
          9828 => x"20253034",
          9829 => x"582d0000",
          9830 => x"25303858",
          9831 => x"20253038",
          9832 => x"582d0000",
          9833 => x"45786563",
          9834 => x"7574696e",
          9835 => x"6720636f",
          9836 => x"64652040",
          9837 => x"20253038",
          9838 => x"78202e2e",
          9839 => x"2e0a0000",
          9840 => x"43616c6c",
          9841 => x"696e6720",
          9842 => x"636f6465",
          9843 => x"20402025",
          9844 => x"30387820",
          9845 => x"2e2e2e0a",
          9846 => x"00000000",
          9847 => x"43616c6c",
          9848 => x"20726574",
          9849 => x"75726e65",
          9850 => x"6420636f",
          9851 => x"64652028",
          9852 => x"2564292e",
          9853 => x"0a000000",
          9854 => x"52657374",
          9855 => x"61727469",
          9856 => x"6e672061",
          9857 => x"70706c69",
          9858 => x"63617469",
          9859 => x"6f6e2e2e",
          9860 => x"2e0a0000",
          9861 => x"436f6c64",
          9862 => x"20726562",
          9863 => x"6f6f7469",
          9864 => x"6e672e2e",
          9865 => x"2e0a0000",
          9866 => x"5a505500",
          9867 => x"62696e00",
          9868 => x"25643a5c",
          9869 => x"25735c25",
          9870 => x"732e2573",
          9871 => x"00000000",
          9872 => x"25643a5c",
          9873 => x"25735c25",
          9874 => x"73000000",
          9875 => x"25643a5c",
          9876 => x"25730000",
          9877 => x"42616420",
          9878 => x"636f6d6d",
          9879 => x"616e642e",
          9880 => x"0a000000",
          9881 => x"52756e6e",
          9882 => x"696e672e",
          9883 => x"2e2e0a00",
          9884 => x"456e6162",
          9885 => x"6c696e67",
          9886 => x"20696e74",
          9887 => x"65727275",
          9888 => x"7074732e",
          9889 => x"2e2e0a00",
          9890 => x"25642f25",
          9891 => x"642f2564",
          9892 => x"2025643a",
          9893 => x"25643a25",
          9894 => x"642e2564",
          9895 => x"25640a00",
          9896 => x"536f4320",
          9897 => x"436f6e66",
          9898 => x"69677572",
          9899 => x"6174696f",
          9900 => x"6e000000",
          9901 => x"20286672",
          9902 => x"6f6d2053",
          9903 => x"6f432063",
          9904 => x"6f6e6669",
          9905 => x"67290000",
          9906 => x"3a0a4465",
          9907 => x"76696365",
          9908 => x"7320696d",
          9909 => x"706c656d",
          9910 => x"656e7465",
          9911 => x"643a0a00",
          9912 => x"20202020",
          9913 => x"57422053",
          9914 => x"4452414d",
          9915 => x"20202825",
          9916 => x"3038583a",
          9917 => x"25303858",
          9918 => x"292e0a00",
          9919 => x"20202020",
          9920 => x"53445241",
          9921 => x"4d202020",
          9922 => x"20202825",
          9923 => x"3038583a",
          9924 => x"25303858",
          9925 => x"292e0a00",
          9926 => x"20202020",
          9927 => x"494e534e",
          9928 => x"20425241",
          9929 => x"4d202825",
          9930 => x"3038583a",
          9931 => x"25303858",
          9932 => x"292e0a00",
          9933 => x"20202020",
          9934 => x"4252414d",
          9935 => x"20202020",
          9936 => x"20202825",
          9937 => x"3038583a",
          9938 => x"25303858",
          9939 => x"292e0a00",
          9940 => x"20202020",
          9941 => x"52414d20",
          9942 => x"20202020",
          9943 => x"20202825",
          9944 => x"3038583a",
          9945 => x"25303858",
          9946 => x"292e0a00",
          9947 => x"20202020",
          9948 => x"53442043",
          9949 => x"41524420",
          9950 => x"20202844",
          9951 => x"65766963",
          9952 => x"6573203d",
          9953 => x"25303264",
          9954 => x"292e0a00",
          9955 => x"20202020",
          9956 => x"54494d45",
          9957 => x"52312020",
          9958 => x"20202854",
          9959 => x"696d6572",
          9960 => x"7320203d",
          9961 => x"25303264",
          9962 => x"292e0a00",
          9963 => x"20202020",
          9964 => x"494e5452",
          9965 => x"20435452",
          9966 => x"4c202843",
          9967 => x"68616e6e",
          9968 => x"656c733d",
          9969 => x"25303264",
          9970 => x"292e0a00",
          9971 => x"20202020",
          9972 => x"57495348",
          9973 => x"424f4e45",
          9974 => x"20425553",
          9975 => x"0a000000",
          9976 => x"20202020",
          9977 => x"57422049",
          9978 => x"32430a00",
          9979 => x"20202020",
          9980 => x"494f4354",
          9981 => x"4c0a0000",
          9982 => x"20202020",
          9983 => x"5053320a",
          9984 => x"00000000",
          9985 => x"20202020",
          9986 => x"5350490a",
          9987 => x"00000000",
          9988 => x"41646472",
          9989 => x"65737365",
          9990 => x"733a0a00",
          9991 => x"20202020",
          9992 => x"43505520",
          9993 => x"52657365",
          9994 => x"74205665",
          9995 => x"63746f72",
          9996 => x"20416464",
          9997 => x"72657373",
          9998 => x"203d2025",
          9999 => x"3038580a",
         10000 => x"00000000",
         10001 => x"20202020",
         10002 => x"43505520",
         10003 => x"4d656d6f",
         10004 => x"72792053",
         10005 => x"74617274",
         10006 => x"20416464",
         10007 => x"72657373",
         10008 => x"203d2025",
         10009 => x"3038580a",
         10010 => x"00000000",
         10011 => x"20202020",
         10012 => x"53746163",
         10013 => x"6b205374",
         10014 => x"61727420",
         10015 => x"41646472",
         10016 => x"65737320",
         10017 => x"20202020",
         10018 => x"203d2025",
         10019 => x"3038580a",
         10020 => x"00000000",
         10021 => x"4d697363",
         10022 => x"3a0a0000",
         10023 => x"20202020",
         10024 => x"5a505520",
         10025 => x"49642020",
         10026 => x"20202020",
         10027 => x"20202020",
         10028 => x"20202020",
         10029 => x"20202020",
         10030 => x"203d2025",
         10031 => x"3034580a",
         10032 => x"00000000",
         10033 => x"20202020",
         10034 => x"53797374",
         10035 => x"656d2043",
         10036 => x"6c6f636b",
         10037 => x"20467265",
         10038 => x"71202020",
         10039 => x"20202020",
         10040 => x"203d2025",
         10041 => x"642e2530",
         10042 => x"34644d48",
         10043 => x"7a0a0000",
         10044 => x"20202020",
         10045 => x"53445241",
         10046 => x"4d20436c",
         10047 => x"6f636b20",
         10048 => x"46726571",
         10049 => x"20202020",
         10050 => x"20202020",
         10051 => x"203d2025",
         10052 => x"642e2530",
         10053 => x"34644d48",
         10054 => x"7a0a0000",
         10055 => x"20202020",
         10056 => x"57697368",
         10057 => x"626f6e65",
         10058 => x"20534452",
         10059 => x"414d2043",
         10060 => x"6c6f636b",
         10061 => x"20467265",
         10062 => x"713d2025",
         10063 => x"642e2530",
         10064 => x"34644d48",
         10065 => x"7a0a0000",
         10066 => x"536d616c",
         10067 => x"6c000000",
         10068 => x"4d656469",
         10069 => x"756d0000",
         10070 => x"466c6578",
         10071 => x"00000000",
         10072 => x"45564f00",
         10073 => x"45564f6d",
         10074 => x"696e0000",
         10075 => x"556e6b6e",
         10076 => x"6f776e00",
         10077 => x"00007ed0",
         10078 => x"01000000",
         10079 => x"00000002",
         10080 => x"00007ecc",
         10081 => x"01000000",
         10082 => x"00000003",
         10083 => x"00007ec8",
         10084 => x"01000000",
         10085 => x"00000004",
         10086 => x"00007ec4",
         10087 => x"01000000",
         10088 => x"00000005",
         10089 => x"00007ec0",
         10090 => x"01000000",
         10091 => x"00000006",
         10092 => x"00007ebc",
         10093 => x"01000000",
         10094 => x"00000007",
         10095 => x"00007eb8",
         10096 => x"01000000",
         10097 => x"00000001",
         10098 => x"00007eb4",
         10099 => x"01000000",
         10100 => x"00000008",
         10101 => x"00007eb0",
         10102 => x"01000000",
         10103 => x"0000000b",
         10104 => x"00007eac",
         10105 => x"01000000",
         10106 => x"00000009",
         10107 => x"00007ea8",
         10108 => x"01000000",
         10109 => x"0000000a",
         10110 => x"00007ea4",
         10111 => x"04000000",
         10112 => x"0000000d",
         10113 => x"00007ea0",
         10114 => x"04000000",
         10115 => x"0000000c",
         10116 => x"00007e9c",
         10117 => x"04000000",
         10118 => x"0000000e",
         10119 => x"00007e98",
         10120 => x"03000000",
         10121 => x"0000000f",
         10122 => x"00007e94",
         10123 => x"04000000",
         10124 => x"0000000f",
         10125 => x"00007e90",
         10126 => x"04000000",
         10127 => x"00000010",
         10128 => x"00007e8c",
         10129 => x"04000000",
         10130 => x"00000011",
         10131 => x"00007e88",
         10132 => x"03000000",
         10133 => x"00000012",
         10134 => x"00007e84",
         10135 => x"03000000",
         10136 => x"00000013",
         10137 => x"00007e80",
         10138 => x"03000000",
         10139 => x"00000014",
         10140 => x"00007e7c",
         10141 => x"03000000",
         10142 => x"00000015",
         10143 => x"1b5b4400",
         10144 => x"1b5b4300",
         10145 => x"1b5b4200",
         10146 => x"1b5b4100",
         10147 => x"1b5b367e",
         10148 => x"1b5b357e",
         10149 => x"1b5b347e",
         10150 => x"1b304600",
         10151 => x"1b5b337e",
         10152 => x"1b5b327e",
         10153 => x"1b5b317e",
         10154 => x"10000000",
         10155 => x"0e000000",
         10156 => x"0d000000",
         10157 => x"0b000000",
         10158 => x"08000000",
         10159 => x"06000000",
         10160 => x"05000000",
         10161 => x"04000000",
         10162 => x"03000000",
         10163 => x"02000000",
         10164 => x"01000000",
         10165 => x"68697374",
         10166 => x"6f727900",
         10167 => x"68697374",
         10168 => x"00000000",
         10169 => x"21000000",
         10170 => x"25303464",
         10171 => x"20202573",
         10172 => x"0a000000",
         10173 => x"4661696c",
         10174 => x"65642074",
         10175 => x"6f207265",
         10176 => x"73657420",
         10177 => x"74686520",
         10178 => x"68697374",
         10179 => x"6f727920",
         10180 => x"66696c65",
         10181 => x"20746f20",
         10182 => x"454f462e",
         10183 => x"0a000000",
         10184 => x"43616e6e",
         10185 => x"6f74206f",
         10186 => x"70656e2f",
         10187 => x"63726561",
         10188 => x"74652068",
         10189 => x"6973746f",
         10190 => x"72792066",
         10191 => x"696c652c",
         10192 => x"20646973",
         10193 => x"61626c69",
         10194 => x"6e672e0a",
         10195 => x"00000000",
         10196 => x"53440000",
         10197 => x"222a2b2c",
         10198 => x"3a3b3c3d",
         10199 => x"3e3f5b5d",
         10200 => x"7c7f0000",
         10201 => x"46415400",
         10202 => x"46415433",
         10203 => x"32000000",
         10204 => x"ebfe904d",
         10205 => x"53444f53",
         10206 => x"352e3000",
         10207 => x"4e4f204e",
         10208 => x"414d4520",
         10209 => x"20202046",
         10210 => x"41543332",
         10211 => x"20202000",
         10212 => x"4e4f204e",
         10213 => x"414d4520",
         10214 => x"20202046",
         10215 => x"41542020",
         10216 => x"20202000",
         10217 => x"00007f50",
         10218 => x"00000000",
         10219 => x"00000000",
         10220 => x"00000000",
         10221 => x"809a4541",
         10222 => x"8e418f80",
         10223 => x"45454549",
         10224 => x"49498e8f",
         10225 => x"9092924f",
         10226 => x"994f5555",
         10227 => x"59999a9b",
         10228 => x"9c9d9e9f",
         10229 => x"41494f55",
         10230 => x"a5a5a6a7",
         10231 => x"a8a9aaab",
         10232 => x"acadaeaf",
         10233 => x"b0b1b2b3",
         10234 => x"b4b5b6b7",
         10235 => x"b8b9babb",
         10236 => x"bcbdbebf",
         10237 => x"c0c1c2c3",
         10238 => x"c4c5c6c7",
         10239 => x"c8c9cacb",
         10240 => x"cccdcecf",
         10241 => x"d0d1d2d3",
         10242 => x"d4d5d6d7",
         10243 => x"d8d9dadb",
         10244 => x"dcdddedf",
         10245 => x"e0e1e2e3",
         10246 => x"e4e5e6e7",
         10247 => x"e8e9eaeb",
         10248 => x"ecedeeef",
         10249 => x"f0f1f2f3",
         10250 => x"f4f5f6f7",
         10251 => x"f8f9fafb",
         10252 => x"fcfdfeff",
         10253 => x"2b2e2c3b",
         10254 => x"3d5b5d2f",
         10255 => x"5c222a3a",
         10256 => x"3c3e3f7c",
         10257 => x"7f000000",
         10258 => x"00010004",
         10259 => x"00100040",
         10260 => x"01000200",
         10261 => x"00000000",
         10262 => x"00010002",
         10263 => x"00040008",
         10264 => x"00100020",
         10265 => x"00000000",
         10266 => x"00000000",
         10267 => x"000074c8",
         10268 => x"01020100",
         10269 => x"00000000",
         10270 => x"00000000",
         10271 => x"000074d0",
         10272 => x"01040100",
         10273 => x"00000000",
         10274 => x"00000000",
         10275 => x"000074d8",
         10276 => x"01140300",
         10277 => x"00000000",
         10278 => x"00000000",
         10279 => x"000074e0",
         10280 => x"012b0300",
         10281 => x"00000000",
         10282 => x"00000000",
         10283 => x"000074e8",
         10284 => x"01300300",
         10285 => x"00000000",
         10286 => x"00000000",
         10287 => x"000074f0",
         10288 => x"013c0400",
         10289 => x"00000000",
         10290 => x"00000000",
         10291 => x"000074f8",
         10292 => x"013d0400",
         10293 => x"00000000",
         10294 => x"00000000",
         10295 => x"00007500",
         10296 => x"013f0400",
         10297 => x"00000000",
         10298 => x"00000000",
         10299 => x"00007508",
         10300 => x"01400400",
         10301 => x"00000000",
         10302 => x"00000000",
         10303 => x"00007510",
         10304 => x"01410400",
         10305 => x"00000000",
         10306 => x"00000000",
         10307 => x"00007514",
         10308 => x"01420400",
         10309 => x"00000000",
         10310 => x"00000000",
         10311 => x"00007518",
         10312 => x"01430400",
         10313 => x"00000000",
         10314 => x"00000000",
         10315 => x"0000751c",
         10316 => x"01500500",
         10317 => x"00000000",
         10318 => x"00000000",
         10319 => x"00007520",
         10320 => x"01510500",
         10321 => x"00000000",
         10322 => x"00000000",
         10323 => x"00007524",
         10324 => x"01540500",
         10325 => x"00000000",
         10326 => x"00000000",
         10327 => x"00007528",
         10328 => x"01550500",
         10329 => x"00000000",
         10330 => x"00000000",
         10331 => x"0000752c",
         10332 => x"01790700",
         10333 => x"00000000",
         10334 => x"00000000",
         10335 => x"00007534",
         10336 => x"01780700",
         10337 => x"00000000",
         10338 => x"00000000",
         10339 => x"00007538",
         10340 => x"01820800",
         10341 => x"00000000",
         10342 => x"00000000",
         10343 => x"00007540",
         10344 => x"01830800",
         10345 => x"00000000",
         10346 => x"00000000",
         10347 => x"00007548",
         10348 => x"01850800",
         10349 => x"00000000",
         10350 => x"00000000",
         10351 => x"00007550",
         10352 => x"01870800",
         10353 => x"00000000",
         10354 => x"00000000",
         10355 => x"00007558",
         10356 => x"018c0900",
         10357 => x"00000000",
         10358 => x"00000000",
         10359 => x"00007560",
         10360 => x"018d0900",
         10361 => x"00000000",
         10362 => x"00000000",
         10363 => x"00007568",
         10364 => x"018e0900",
         10365 => x"00000000",
         10366 => x"00000000",
         10367 => x"00007570",
         10368 => x"018f0900",
         10369 => x"00000000",
         10370 => x"00000000",
         10371 => x"00000000",
         10372 => x"00000000",
         10373 => x"00007fff",
         10374 => x"00000000",
         10375 => x"00007fff",
         10376 => x"00010000",
         10377 => x"00007fff",
         10378 => x"00010000",
         10379 => x"00810000",
         10380 => x"01000000",
         10381 => x"017fffff",
         10382 => x"00000000",
         10383 => x"00000000",
         10384 => x"00007800",
         10385 => x"00000000",
         10386 => x"05f5e100",
         10387 => x"05f5e100",
         10388 => x"05f5e100",
         10389 => x"00000000",
         10390 => x"01010101",
         10391 => x"01010101",
         10392 => x"01011001",
         10393 => x"01000000",
         10394 => x"00000000",
         10395 => x"00000000",
         10396 => x"00000000",
         10397 => x"00000000",
         10398 => x"00000000",
         10399 => x"00000000",
         10400 => x"00000000",
         10401 => x"00000000",
         10402 => x"00000000",
         10403 => x"00000000",
         10404 => x"00000000",
         10405 => x"00000000",
         10406 => x"00000000",
         10407 => x"00000000",
         10408 => x"00000000",
         10409 => x"00000000",
         10410 => x"00000000",
         10411 => x"00000000",
         10412 => x"00000000",
         10413 => x"00000000",
         10414 => x"00000000",
         10415 => x"00000000",
         10416 => x"00000000",
         10417 => x"00000000",
         10418 => x"00007ed4",
         10419 => x"01000000",
         10420 => x"00007edc",
         10421 => x"01000000",
         10422 => x"00007ee4",
         10423 => x"02000000",
         10424 => x"00000000",
         10425 => x"00000000",
         10426 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

